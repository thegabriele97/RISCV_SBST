
library IEEE;
library c6288;

use IEEE.std_logic_1164.all;
use c6288.gate_lib.all;

entity c6288 is

   port( datai : in std_logic_vector(31 downto 0);
         datao : out std_logic_vector(31 downto 0));
         
end c6288;

architecture SYN_USE_DEFA_ARCH_NAME of c6288 is

signal   G_1GAT, G_18GAT, G_35GAT, G_52GAT, G_69GAT, G_86GAT, G_103GAT, 
         G_120GAT, G_137GAT, G_154GAT, G_171GAT, G_188GAT, G_205GAT, G_222GAT, 
         G_239GAT, G_256GAT, G_273GAT, G_290GAT, G_307GAT, G_324GAT, G_341GAT, 
         G_358GAT, G_375GAT, G_392GAT, G_409GAT, G_426GAT, G_443GAT, G_460GAT, 
         G_477GAT, G_494GAT, G_511GAT, G_528GAT : std_logic;
signal   G_545GAT_PO, G_1581GAT_PO, G_1901GAT_PO, G_2223GAT_PO, G_2548GAT_PO, G_2877GAT_PO, 
         G_3211GAT_PO, G_3552GAT_PO, G_3895GAT_PO, G_4241GAT_PO, G_4591GAT_PO, 
         G_4946GAT_PO, G_5308GAT_PO, G_5672GAT_PO, G_5971GAT_PO, G_6123GAT_PO, 
         G_6150GAT_PO, G_6160GAT_PO, G_6170GAT_PO, G_6180GAT_PO, G_6190GAT_PO, 
         G_6200GAT_PO, G_6210GAT_PO, G_6220GAT_PO, G_6230GAT_PO, G_6240GAT_PO, 
         G_6250GAT_PO, G_6260GAT_PO, G_6270GAT_PO, G_6280GAT_PO, G_6287GAT_PO, 
         G_6288GAT_PO : std_logic;









   component Nor_gate
      port( I1, I2 : in std_logic;  O : out std_logic);
   end component;
   
   component Inv_gate
      port( I1 : in std_logic;  O : out std_logic);
   end component;
   
   component And_gate
      port( I1, I2 : in std_logic;  O : out std_logic);
   end component;
   
   signal G_6286GAT_OUT, G_6285GAT_OUT, G_6281GAT_OUT, G_6277GAT_OUT, 
      G_6276GAT_OUT, G_6275GAT_OUT, G_6271GAT_OUT, G_6267GAT_OUT, G_6266GAT_OUT
      , G_6265GAT_OUT, G_6261GAT_OUT, G_6257GAT_OUT, G_6256GAT_OUT, 
      G_6255GAT_OUT, G_6251GAT_OUT, G_6247GAT_OUT, G_6246GAT_OUT, G_6245GAT_OUT
      , G_6241GAT_OUT, G_6237GAT_OUT, G_6236GAT_OUT, G_6235GAT_OUT, 
      G_6231GAT_OUT, G_6227GAT_OUT, G_6226GAT_OUT, G_6225GAT_OUT, G_6221GAT_OUT
      , G_6217GAT_OUT, G_6216GAT_OUT, G_6215GAT_OUT, G_6211GAT_OUT, 
      G_6207GAT_OUT, G_6206GAT_OUT, G_6205GAT_OUT, G_6201GAT_OUT, G_6197GAT_OUT
      , G_6196GAT_OUT, G_6195GAT_OUT, G_6191GAT_OUT, G_6187GAT_OUT, 
      G_6186GAT_OUT, G_6185GAT_OUT, G_6181GAT_OUT, G_6177GAT_OUT, G_6176GAT_OUT
      , G_6175GAT_OUT, G_6171GAT_OUT, G_6167GAT_OUT, G_6166GAT_OUT, 
      G_6165GAT_OUT, G_6161GAT_OUT, G_6157GAT_OUT, G_6156GAT_OUT, G_6155GAT_OUT
      , G_6151GAT_OUT, G_6147GAT_OUT, G_6146GAT_OUT, G_6145GAT_OUT, 
      G_6141GAT_OUT, G_6138GAT_OUT, G_6135GAT_OUT, G_6134GAT_OUT, G_6133GAT_OUT
      , G_6130GAT_OUT, G_6129GAT_OUT, G_6128GAT_OUT, G_6124GAT_OUT, 
      G_6120GAT_OUT, G_6119GAT_OUT, G_6118GAT_OUT, G_6114GAT_OUT, G_6111GAT_OUT
      , G_6108GAT_OUT, G_6107GAT_OUT, G_6106GAT_OUT, G_6103GAT_OUT, 
      G_6102GAT_OUT, G_6101GAT_OUT, G_6097GAT_OUT, G_6094GAT_OUT, G_6091GAT_OUT
      , G_6090GAT_OUT, G_6089GAT_OUT, G_6085GAT_OUT, G_6082GAT_OUT, 
      G_6081GAT_OUT, G_6080GAT_OUT, G_6076GAT_OUT, G_6073GAT_OUT, G_6070GAT_OUT
      , G_6069GAT_OUT, G_6068GAT_OUT, G_6064GAT_OUT, G_6061GAT_OUT, 
      G_6058GAT_OUT, G_6057GAT_OUT, G_6056GAT_OUT, G_6052GAT_OUT, G_6049GAT_OUT
      , G_6046GAT_OUT, G_6045GAT_OUT, G_6044GAT_OUT, G_6040GAT_OUT, 
      G_6037GAT_OUT, G_6036GAT_OUT, G_6035GAT_OUT, G_6032GAT_OUT, G_6031GAT_OUT
      , G_6030GAT_OUT, G_6026GAT_OUT, G_6023GAT_OUT, G_6020GAT_OUT, 
      G_6019GAT_OUT, G_6018GAT_OUT, G_6014GAT_OUT, G_6011GAT_OUT, G_6010GAT_OUT
      , G_6009GAT_OUT, G_6005GAT_OUT, G_6002GAT_OUT, G_6001GAT_OUT, 
      G_6000GAT_OUT, G_5996GAT_OUT, G_5993GAT_OUT, G_5990GAT_OUT, G_5989GAT_OUT
      , G_5988GAT_OUT, G_5984GAT_OUT, G_5981GAT_OUT, G_5980GAT_OUT, 
      G_5979GAT_OUT, G_5975GAT_OUT, G_5972GAT_OUT, G_5968GAT_OUT, G_5967GAT_OUT
      , G_5966GAT_OUT, G_5962GAT_OUT, G_5959GAT_OUT, G_5956GAT_OUT, 
      G_5955GAT_OUT, G_5954GAT_OUT, G_5950GAT_OUT, G_5947GAT_OUT, G_5946GAT_OUT
      , G_5945GAT_OUT, G_5941GAT_OUT, G_5938GAT_OUT, G_5935GAT_OUT, 
      G_5934GAT_OUT, G_5933GAT_OUT, G_5930GAT_OUT, G_5929GAT_OUT, G_5928GAT_OUT
      , G_5925GAT_OUT, G_5924GAT_OUT, G_5923GAT_OUT, G_5919GAT_OUT, 
      G_5916GAT_OUT, G_5913GAT_OUT, G_5912GAT_OUT, G_5911GAT_OUT, G_5907GAT_OUT
      , G_5904GAT_OUT, G_5903GAT_OUT, G_5902GAT_OUT, G_5898GAT_OUT, 
      G_5895GAT_OUT, G_5892GAT_OUT, G_5891GAT_OUT, G_5890GAT_OUT, G_5886GAT_OUT
      , G_5882GAT_OUT, G_5879GAT_OUT, G_5878GAT_OUT, G_5877GAT_OUT, 
      G_5873GAT_OUT, G_5870GAT_OUT, G_5867GAT_OUT, G_5866GAT_OUT, G_5865GAT_OUT
      , G_5861GAT_OUT, G_5858GAT_OUT, G_5857GAT_OUT, G_5856GAT_OUT, 
      G_5852GAT_OUT, G_5849GAT_OUT, G_5846GAT_OUT, G_5845GAT_OUT, G_5844GAT_OUT
      , G_5840GAT_OUT, G_5837GAT_OUT, G_5834GAT_OUT, G_5831GAT_OUT, 
      G_5830GAT_OUT, G_5829GAT_OUT, G_5825GAT_OUT, G_5822GAT_OUT, G_5819GAT_OUT
      , G_5818GAT_OUT, G_5817GAT_OUT, G_5813GAT_OUT, G_5810GAT_OUT, 
      G_5809GAT_OUT, G_5808GAT_OUT, G_5804GAT_OUT, G_5801GAT_OUT, G_5798GAT_OUT
      , G_5797GAT_OUT, G_5796GAT_OUT, G_5792GAT_OUT, G_5789GAT_OUT, 
      G_5788GAT_OUT, G_5787GAT_OUT, G_5786GAT_OUT, G_5785GAT_OUT, G_5782GAT_OUT
      , G_5781GAT_OUT, G_5780GAT_OUT, G_5776GAT_OUT, G_5773GAT_OUT, 
      G_5770GAT_OUT, G_5769GAT_OUT, G_5768GAT_OUT, G_5764GAT_OUT, G_5761GAT_OUT
      , G_5760GAT_OUT, G_5759GAT_OUT, G_5755GAT_OUT, G_5752GAT_OUT, 
      G_5749GAT_OUT, G_5748GAT_OUT, G_5747GAT_OUT, G_5743GAT_OUT, G_5740GAT_OUT
      , G_5739GAT_OUT, G_5738GAT_OUT, G_5734GAT_OUT, G_5730GAT_OUT, 
      G_5727GAT_OUT, G_5726GAT_OUT, G_5725GAT_OUT, G_5721GAT_OUT, G_5718GAT_OUT
      , G_5715GAT_OUT, G_5714GAT_OUT, G_5713GAT_OUT, G_5709GAT_OUT, 
      G_5706GAT_OUT, G_5705GAT_OUT, G_5704GAT_OUT, G_5700GAT_OUT, G_5697GAT_OUT
      , G_5694GAT_OUT, G_5693GAT_OUT, G_5692GAT_OUT, G_5688GAT_OUT, 
      G_5685GAT_OUT, G_5684GAT_OUT, G_5683GAT_OUT, G_5679GAT_OUT, G_5676GAT_OUT
      , G_5673GAT_OUT, G_5671GAT_OUT, G_5670GAT_OUT, G_5666GAT_OUT, 
      G_5663GAT_OUT, G_5660GAT_OUT, G_5659GAT_OUT, G_5658GAT_OUT, G_5654GAT_OUT
      , G_5651GAT_OUT, G_5650GAT_OUT, G_5649GAT_OUT, G_5645GAT_OUT, 
      G_5642GAT_OUT, G_5639GAT_OUT, G_5638GAT_OUT, G_5637GAT_OUT, G_5633GAT_OUT
      , G_5630GAT_OUT, G_5629GAT_OUT, G_5628GAT_OUT, G_5624GAT_OUT, 
      G_5621GAT_OUT, G_5618GAT_OUT, G_5617GAT_OUT, G_5616GAT_OUT, G_5613GAT_OUT
      , G_5612GAT_OUT, G_5611GAT_OUT, G_5608GAT_OUT, G_5607GAT_OUT, 
      G_5606GAT_OUT, G_5602GAT_OUT, G_5599GAT_OUT, G_5596GAT_OUT, G_5595GAT_OUT
      , G_5594GAT_OUT, G_5590GAT_OUT, G_5587GAT_OUT, G_5586GAT_OUT, 
      G_5585GAT_OUT, G_5581GAT_OUT, G_5578GAT_OUT, G_5575GAT_OUT, G_5574GAT_OUT
      , G_5573GAT_OUT, G_5569GAT_OUT, G_5566GAT_OUT, G_5565GAT_OUT, 
      G_5564GAT_OUT, G_5560GAT_OUT, G_5557GAT_OUT, G_5554GAT_OUT, G_5553GAT_OUT
      , G_5552GAT_OUT, G_5548GAT_OUT, G_5544GAT_OUT, G_5540GAT_OUT, 
      G_5537GAT_OUT, G_5536GAT_OUT, G_5535GAT_OUT, G_5531GAT_OUT, G_5528GAT_OUT
      , G_5527GAT_OUT, G_5526GAT_OUT, G_5522GAT_OUT, G_5519GAT_OUT, 
      G_5516GAT_OUT, G_5515GAT_OUT, G_5514GAT_OUT, G_5510GAT_OUT, G_5507GAT_OUT
      , G_5506GAT_OUT, G_5505GAT_OUT, G_5501GAT_OUT, G_5498GAT_OUT, 
      G_5495GAT_OUT, G_5494GAT_OUT, G_5493GAT_OUT, G_5489GAT_OUT, G_5486GAT_OUT
      , G_5483GAT_OUT, G_5480GAT_OUT, G_5476GAT_OUT, G_5473GAT_OUT, 
      G_5472GAT_OUT, G_5471GAT_OUT, G_5467GAT_OUT, G_5464GAT_OUT, G_5461GAT_OUT
      , G_5460GAT_OUT, G_5459GAT_OUT, G_5455GAT_OUT, G_5452GAT_OUT, 
      G_5451GAT_OUT, G_5450GAT_OUT, G_5446GAT_OUT, G_5443GAT_OUT, G_5440GAT_OUT
      , G_5439GAT_OUT, G_5438GAT_OUT, G_5434GAT_OUT, G_5431GAT_OUT, 
      G_5430GAT_OUT, G_5429GAT_OUT, G_5428GAT_OUT, G_5427GAT_OUT, G_5426GAT_OUT
      , G_5425GAT_OUT, G_5422GAT_OUT, G_5421GAT_OUT, G_5420GAT_OUT, 
      G_5416GAT_OUT, G_5413GAT_OUT, G_5410GAT_OUT, G_5409GAT_OUT, G_5408GAT_OUT
      , G_5404GAT_OUT, G_5401GAT_OUT, G_5400GAT_OUT, G_5399GAT_OUT, 
      G_5395GAT_OUT, G_5392GAT_OUT, G_5389GAT_OUT, G_5388GAT_OUT, G_5387GAT_OUT
      , G_5383GAT_OUT, G_5380GAT_OUT, G_5379GAT_OUT, G_5378GAT_OUT, 
      G_5374GAT_OUT, G_5370GAT_OUT, G_5366GAT_OUT, G_5365GAT_OUT, G_5364GAT_OUT
      , G_5360GAT_OUT, G_5357GAT_OUT, G_5354GAT_OUT, G_5353GAT_OUT, 
      G_5352GAT_OUT, G_5348GAT_OUT, G_5345GAT_OUT, G_5344GAT_OUT, G_5343GAT_OUT
      , G_5339GAT_OUT, G_5336GAT_OUT, G_5333GAT_OUT, G_5332GAT_OUT, 
      G_5331GAT_OUT, G_5327GAT_OUT, G_5324GAT_OUT, G_5323GAT_OUT, G_5322GAT_OUT
      , G_5318GAT_OUT, G_5315GAT_OUT, G_5312GAT_OUT, G_5309GAT_OUT, 
      G_5304GAT_OUT, G_5301GAT_OUT, G_5298GAT_OUT, G_5297GAT_OUT, G_5296GAT_OUT
      , G_5292GAT_OUT, G_5289GAT_OUT, G_5288GAT_OUT, G_5287GAT_OUT, 
      G_5283GAT_OUT, G_5280GAT_OUT, G_5277GAT_OUT, G_5276GAT_OUT, G_5275GAT_OUT
      , G_5271GAT_OUT, G_5268GAT_OUT, G_5267GAT_OUT, G_5266GAT_OUT, 
      G_5262GAT_OUT, G_5259GAT_OUT, G_5256GAT_OUT, G_5255GAT_OUT, G_5254GAT_OUT
      , G_5251GAT_OUT, G_5250GAT_OUT, G_5249GAT_OUT, G_5246GAT_OUT, 
      G_5245GAT_OUT, G_5244GAT_OUT, G_5241GAT_OUT, G_5240GAT_OUT, G_5239GAT_OUT
      , G_5236GAT_OUT, G_5235GAT_OUT, G_5234GAT_OUT, G_5230GAT_OUT, 
      G_5227GAT_OUT, G_5226GAT_OUT, G_5225GAT_OUT, G_5221GAT_OUT, G_5218GAT_OUT
      , G_5215GAT_OUT, G_5214GAT_OUT, G_5213GAT_OUT, G_5209GAT_OUT, 
      G_5206GAT_OUT, G_5205GAT_OUT, G_5204GAT_OUT, G_5200GAT_OUT, G_5197GAT_OUT
      , G_5194GAT_OUT, G_5193GAT_OUT, G_5192GAT_OUT, G_5188GAT_OUT, 
      G_5184GAT_OUT, G_5180GAT_OUT, G_5176GAT_OUT, G_5172GAT_OUT, G_5169GAT_OUT
      , G_5168GAT_OUT, G_5167GAT_OUT, G_5163GAT_OUT, G_5160GAT_OUT, 
      G_5157GAT_OUT, G_5156GAT_OUT, G_5155GAT_OUT, G_5151GAT_OUT, G_5148GAT_OUT
      , G_5147GAT_OUT, G_5146GAT_OUT, G_5142GAT_OUT, G_5139GAT_OUT, 
      G_5136GAT_OUT, G_5135GAT_OUT, G_5134GAT_OUT, G_5130GAT_OUT, G_5127GAT_OUT
      , G_5124GAT_OUT, G_5121GAT_OUT, G_5118GAT_OUT, G_5115GAT_OUT, 
      G_5114GAT_OUT, G_5113GAT_OUT, G_5109GAT_OUT, G_5106GAT_OUT, G_5103GAT_OUT
      , G_5102GAT_OUT, G_5101GAT_OUT, G_5097GAT_OUT, G_5094GAT_OUT, 
      G_5093GAT_OUT, G_5092GAT_OUT, G_5088GAT_OUT, G_5085GAT_OUT, G_5082GAT_OUT
      , G_5081GAT_OUT, G_5080GAT_OUT, G_5076GAT_OUT, G_5073GAT_OUT, 
      G_5072GAT_OUT, G_5071GAT_OUT, G_5070GAT_OUT, G_5069GAT_OUT, G_5068GAT_OUT
      , G_5067GAT_OUT, G_5066GAT_OUT, G_5065GAT_OUT, G_5064GAT_OUT, 
      G_5063GAT_OUT, G_5059GAT_OUT, G_5056GAT_OUT, G_5053GAT_OUT, G_5052GAT_OUT
      , G_5051GAT_OUT, G_5047GAT_OUT, G_5044GAT_OUT, G_5043GAT_OUT, 
      G_5042GAT_OUT, G_5038GAT_OUT, G_5035GAT_OUT, G_5032GAT_OUT, G_5031GAT_OUT
      , G_5030GAT_OUT, G_5026GAT_OUT, G_5023GAT_OUT, G_5022GAT_OUT, 
      G_5021GAT_OUT, G_5017GAT_OUT, G_5013GAT_OUT, G_5009GAT_OUT, G_5005GAT_OUT
      , G_5001GAT_OUT, G_4998GAT_OUT, G_4995GAT_OUT, G_4994GAT_OUT, 
      G_4993GAT_OUT, G_4989GAT_OUT, G_4986GAT_OUT, G_4985GAT_OUT, G_4984GAT_OUT
      , G_4980GAT_OUT, G_4977GAT_OUT, G_4974GAT_OUT, G_4973GAT_OUT, 
      G_4972GAT_OUT, G_4968GAT_OUT, G_4965GAT_OUT, G_4964GAT_OUT, G_4963GAT_OUT
      , G_4959GAT_OUT, G_4956GAT_OUT, G_4953GAT_OUT, G_4950GAT_OUT, 
      G_4947GAT_OUT, G_4943GAT_OUT, G_4942GAT_OUT, G_4941GAT_OUT, G_4937GAT_OUT
      , G_4934GAT_OUT, G_4933GAT_OUT, G_4932GAT_OUT, G_4928GAT_OUT, 
      G_4925GAT_OUT, G_4922GAT_OUT, G_4921GAT_OUT, G_4920GAT_OUT, G_4916GAT_OUT
      , G_4913GAT_OUT, G_4912GAT_OUT, G_4911GAT_OUT, G_4907GAT_OUT, 
      G_4904GAT_OUT, G_4901GAT_OUT, G_4900GAT_OUT, G_4899GAT_OUT, G_4896GAT_OUT
      , G_4895GAT_OUT, G_4894GAT_OUT, G_4891GAT_OUT, G_4890GAT_OUT, 
      G_4889GAT_OUT, G_4886GAT_OUT, G_4885GAT_OUT, G_4884GAT_OUT, G_4881GAT_OUT
      , G_4880GAT_OUT, G_4879GAT_OUT, G_4875GAT_OUT, G_4872GAT_OUT, 
      G_4871GAT_OUT, G_4870GAT_OUT, G_4866GAT_OUT, G_4863GAT_OUT, G_4860GAT_OUT
      , G_4859GAT_OUT, G_4858GAT_OUT, G_4854GAT_OUT, G_4851GAT_OUT, 
      G_4850GAT_OUT, G_4849GAT_OUT, G_4845GAT_OUT, G_4842GAT_OUT, G_4839GAT_OUT
      , G_4838GAT_OUT, G_4837GAT_OUT, G_4833GAT_OUT, G_4829GAT_OUT, 
      G_4825GAT_OUT, G_4821GAT_OUT, G_4817GAT_OUT, G_4814GAT_OUT, G_4813GAT_OUT
      , G_4812GAT_OUT, G_4808GAT_OUT, G_4805GAT_OUT, G_4802GAT_OUT, 
      G_4801GAT_OUT, G_4800GAT_OUT, G_4796GAT_OUT, G_4793GAT_OUT, G_4792GAT_OUT
      , G_4791GAT_OUT, G_4787GAT_OUT, G_4784GAT_OUT, G_4781GAT_OUT, 
      G_4780GAT_OUT, G_4779GAT_OUT, G_4775GAT_OUT, G_4772GAT_OUT, G_4769GAT_OUT
      , G_4766GAT_OUT, G_4763GAT_OUT, G_4760GAT_OUT, G_4759GAT_OUT, 
      G_4758GAT_OUT, G_4754GAT_OUT, G_4751GAT_OUT, G_4748GAT_OUT, G_4747GAT_OUT
      , G_4746GAT_OUT, G_4742GAT_OUT, G_4739GAT_OUT, G_4738GAT_OUT, 
      G_4737GAT_OUT, G_4733GAT_OUT, G_4730GAT_OUT, G_4727GAT_OUT, G_4726GAT_OUT
      , G_4725GAT_OUT, G_4721GAT_OUT, G_4718GAT_OUT, G_4717GAT_OUT, 
      G_4716GAT_OUT, G_4715GAT_OUT, G_4714GAT_OUT, G_4713GAT_OUT, G_4712GAT_OUT
      , G_4711GAT_OUT, G_4710GAT_OUT, G_4709GAT_OUT, G_4708GAT_OUT, 
      G_4704GAT_OUT, G_4701GAT_OUT, G_4698GAT_OUT, G_4697GAT_OUT, G_4696GAT_OUT
      , G_4692GAT_OUT, G_4689GAT_OUT, G_4688GAT_OUT, G_4687GAT_OUT, 
      G_4683GAT_OUT, G_4680GAT_OUT, G_4677GAT_OUT, G_4676GAT_OUT, G_4675GAT_OUT
      , G_4671GAT_OUT, G_4668GAT_OUT, G_4667GAT_OUT, G_4666GAT_OUT, 
      G_4662GAT_OUT, G_4658GAT_OUT, G_4654GAT_OUT, G_4650GAT_OUT, G_4646GAT_OUT
      , G_4643GAT_OUT, G_4642GAT_OUT, G_4641GAT_OUT, G_4637GAT_OUT, 
      G_4634GAT_OUT, G_4633GAT_OUT, G_4632GAT_OUT, G_4628GAT_OUT, G_4625GAT_OUT
      , G_4622GAT_OUT, G_4621GAT_OUT, G_4620GAT_OUT, G_4616GAT_OUT, 
      G_4613GAT_OUT, G_4612GAT_OUT, G_4611GAT_OUT, G_4607GAT_OUT, G_4604GAT_OUT
      , G_4601GAT_OUT, G_4598GAT_OUT, G_4595GAT_OUT, G_4592GAT_OUT, 
      G_4587GAT_OUT, G_4584GAT_OUT, G_4583GAT_OUT, G_4582GAT_OUT, G_4578GAT_OUT
      , G_4575GAT_OUT, G_4572GAT_OUT, G_4571GAT_OUT, G_4570GAT_OUT, 
      G_4566GAT_OUT, G_4563GAT_OUT, G_4562GAT_OUT, G_4561GAT_OUT, G_4557GAT_OUT
      , G_4554GAT_OUT, G_4551GAT_OUT, G_4550GAT_OUT, G_4549GAT_OUT, 
      G_4546GAT_OUT, G_4545GAT_OUT, G_4544GAT_OUT, G_4541GAT_OUT, G_4540GAT_OUT
      , G_4539GAT_OUT, G_4536GAT_OUT, G_4535GAT_OUT, G_4534GAT_OUT, 
      G_4531GAT_OUT, G_4530GAT_OUT, G_4529GAT_OUT, G_4526GAT_OUT, G_4525GAT_OUT
      , G_4524GAT_OUT, G_4521GAT_OUT, G_4520GAT_OUT, G_4519GAT_OUT, 
      G_4515GAT_OUT, G_4512GAT_OUT, G_4509GAT_OUT, G_4508GAT_OUT, G_4507GAT_OUT
      , G_4503GAT_OUT, G_4500GAT_OUT, G_4499GAT_OUT, G_4498GAT_OUT, 
      G_4494GAT_OUT, G_4491GAT_OUT, G_4488GAT_OUT, G_4487GAT_OUT, G_4486GAT_OUT
      , G_4482GAT_OUT, G_4478GAT_OUT, G_4474GAT_OUT, G_4470GAT_OUT, 
      G_4466GAT_OUT, G_4462GAT_OUT, G_4461GAT_OUT, G_4460GAT_OUT, G_4456GAT_OUT
      , G_4453GAT_OUT, G_4450GAT_OUT, G_4449GAT_OUT, G_4448GAT_OUT, 
      G_4444GAT_OUT, G_4441GAT_OUT, G_4440GAT_OUT, G_4439GAT_OUT, G_4435GAT_OUT
      , G_4432GAT_OUT, G_4429GAT_OUT, G_4428GAT_OUT, G_4427GAT_OUT, 
      G_4423GAT_OUT, G_4420GAT_OUT, G_4417GAT_OUT, G_4414GAT_OUT, G_4411GAT_OUT
      , G_4408GAT_OUT, G_4405GAT_OUT, G_4401GAT_OUT, G_4398GAT_OUT, 
      G_4395GAT_OUT, G_4394GAT_OUT, G_4393GAT_OUT, G_4389GAT_OUT, G_4386GAT_OUT
      , G_4385GAT_OUT, G_4384GAT_OUT, G_4380GAT_OUT, G_4377GAT_OUT, 
      G_4374GAT_OUT, G_4373GAT_OUT, G_4372GAT_OUT, G_4368GAT_OUT, G_4365GAT_OUT
      , G_4364GAT_OUT, G_4363GAT_OUT, G_4362GAT_OUT, G_4361GAT_OUT, 
      G_4360GAT_OUT, G_4359GAT_OUT, G_4358GAT_OUT, G_4357GAT_OUT, G_4356GAT_OUT
      , G_4355GAT_OUT, G_4354GAT_OUT, G_4353GAT_OUT, G_4350GAT_OUT, 
      G_4349GAT_OUT, G_4348GAT_OUT, G_4344GAT_OUT, G_4341GAT_OUT, G_4340GAT_OUT
      , G_4339GAT_OUT, G_4335GAT_OUT, G_4332GAT_OUT, G_4329GAT_OUT, 
      G_4328GAT_OUT, G_4327GAT_OUT, G_4323GAT_OUT, G_4320GAT_OUT, G_4319GAT_OUT
      , G_4318GAT_OUT, G_4314GAT_OUT, G_4310GAT_OUT, G_4306GAT_OUT, 
      G_4302GAT_OUT, G_4298GAT_OUT, G_4294GAT_OUT, G_4290GAT_OUT, G_4287GAT_OUT
      , G_4286GAT_OUT, G_4285GAT_OUT, G_4281GAT_OUT, G_4278GAT_OUT, 
      G_4275GAT_OUT, G_4274GAT_OUT, G_4273GAT_OUT, G_4269GAT_OUT, G_4266GAT_OUT
      , G_4265GAT_OUT, G_4264GAT_OUT, G_4260GAT_OUT, G_4257GAT_OUT, 
      G_4254GAT_OUT, G_4251GAT_OUT, G_4248GAT_OUT, G_4245GAT_OUT, G_4242GAT_OUT
      , G_4238GAT_OUT, G_4237GAT_OUT, G_4236GAT_OUT, G_4232GAT_OUT, 
      G_4229GAT_OUT, G_4226GAT_OUT, G_4225GAT_OUT, G_4224GAT_OUT, G_4220GAT_OUT
      , G_4217GAT_OUT, G_4216GAT_OUT, G_4215GAT_OUT, G_4211GAT_OUT, 
      G_4208GAT_OUT, G_4205GAT_OUT, G_4204GAT_OUT, G_4203GAT_OUT, G_4200GAT_OUT
      , G_4199GAT_OUT, G_4198GAT_OUT, G_4195GAT_OUT, G_4194GAT_OUT, 
      G_4193GAT_OUT, G_4190GAT_OUT, G_4189GAT_OUT, G_4188GAT_OUT, G_4185GAT_OUT
      , G_4184GAT_OUT, G_4183GAT_OUT, G_4180GAT_OUT, G_4179GAT_OUT, 
      G_4178GAT_OUT, G_4175GAT_OUT, G_4174GAT_OUT, G_4173GAT_OUT, G_4172GAT_OUT
      , G_4171GAT_OUT, G_4167GAT_OUT, G_4164GAT_OUT, G_4161GAT_OUT, 
      G_4160GAT_OUT, G_4159GAT_OUT, G_4155GAT_OUT, G_4152GAT_OUT, G_4151GAT_OUT
      , G_4150GAT_OUT, G_4146GAT_OUT, G_4143GAT_OUT, G_4140GAT_OUT, 
      G_4139GAT_OUT, G_4138GAT_OUT, G_4134GAT_OUT, G_4130GAT_OUT, G_4126GAT_OUT
      , G_4122GAT_OUT, G_4118GAT_OUT, G_4114GAT_OUT, G_4110GAT_OUT, 
      G_4106GAT_OUT, G_4103GAT_OUT, G_4100GAT_OUT, G_4099GAT_OUT, G_4098GAT_OUT
      , G_4094GAT_OUT, G_4091GAT_OUT, G_4090GAT_OUT, G_4089GAT_OUT, 
      G_4085GAT_OUT, G_4082GAT_OUT, G_4079GAT_OUT, G_4078GAT_OUT, G_4077GAT_OUT
      , G_4073GAT_OUT, G_4070GAT_OUT, G_4067GAT_OUT, G_4064GAT_OUT, 
      G_4061GAT_OUT, G_4058GAT_OUT, G_4055GAT_OUT, G_4052GAT_OUT, G_4049GAT_OUT
      , G_4048GAT_OUT, G_4047GAT_OUT, G_4043GAT_OUT, G_4040GAT_OUT, 
      G_4039GAT_OUT, G_4038GAT_OUT, G_4034GAT_OUT, G_4031GAT_OUT, G_4028GAT_OUT
      , G_4027GAT_OUT, G_4026GAT_OUT, G_4022GAT_OUT, G_4019GAT_OUT, 
      G_4018GAT_OUT, G_4017GAT_OUT, G_4016GAT_OUT, G_4015GAT_OUT, G_4014GAT_OUT
      , G_4013GAT_OUT, G_4012GAT_OUT, G_4011GAT_OUT, G_4010GAT_OUT, 
      G_4009GAT_OUT, G_4008GAT_OUT, G_4007GAT_OUT, G_4006GAT_OUT, G_4005GAT_OUT
      , G_4001GAT_OUT, G_3998GAT_OUT, G_3997GAT_OUT, G_3996GAT_OUT, 
      G_3992GAT_OUT, G_3989GAT_OUT, G_3986GAT_OUT, G_3985GAT_OUT, G_3984GAT_OUT
      , G_3980GAT_OUT, G_3977GAT_OUT, G_3976GAT_OUT, G_3975GAT_OUT, 
      G_3971GAT_OUT, G_3967GAT_OUT, G_3963GAT_OUT, G_3959GAT_OUT, G_3955GAT_OUT
      , G_3951GAT_OUT, G_3947GAT_OUT, G_3944GAT_OUT, G_3943GAT_OUT, 
      G_3942GAT_OUT, G_3938GAT_OUT, G_3935GAT_OUT, G_3932GAT_OUT, G_3931GAT_OUT
      , G_3930GAT_OUT, G_3926GAT_OUT, G_3923GAT_OUT, G_3922GAT_OUT, 
      G_3921GAT_OUT, G_3917GAT_OUT, G_3914GAT_OUT, G_3911GAT_OUT, G_3908GAT_OUT
      , G_3905GAT_OUT, G_3902GAT_OUT, G_3899GAT_OUT, G_3896GAT_OUT, 
      G_3894GAT_OUT, G_3893GAT_OUT, G_3889GAT_OUT, G_3886GAT_OUT, G_3883GAT_OUT
      , G_3882GAT_OUT, G_3881GAT_OUT, G_3877GAT_OUT, G_3874GAT_OUT, 
      G_3873GAT_OUT, G_3872GAT_OUT, G_3868GAT_OUT, G_3865GAT_OUT, G_3862GAT_OUT
      , G_3861GAT_OUT, G_3860GAT_OUT, G_3857GAT_OUT, G_3856GAT_OUT, 
      G_3855GAT_OUT, G_3852GAT_OUT, G_3851GAT_OUT, G_3850GAT_OUT, G_3847GAT_OUT
      , G_3846GAT_OUT, G_3845GAT_OUT, G_3842GAT_OUT, G_3841GAT_OUT, 
      G_3840GAT_OUT, G_3837GAT_OUT, G_3836GAT_OUT, G_3835GAT_OUT, G_3832GAT_OUT
      , G_3831GAT_OUT, G_3830GAT_OUT, G_3827GAT_OUT, G_3826GAT_OUT, 
      G_3825GAT_OUT, G_3821GAT_OUT, G_3818GAT_OUT, G_3815GAT_OUT, G_3814GAT_OUT
      , G_3813GAT_OUT, G_3809GAT_OUT, G_3806GAT_OUT, G_3805GAT_OUT, 
      G_3804GAT_OUT, G_3800GAT_OUT, G_3797GAT_OUT, G_3794GAT_OUT, G_3793GAT_OUT
      , G_3792GAT_OUT, G_3788GAT_OUT, G_3784GAT_OUT, G_3780GAT_OUT, 
      G_3776GAT_OUT, G_3772GAT_OUT, G_3768GAT_OUT, G_3764GAT_OUT, G_3760GAT_OUT
      , G_3757GAT_OUT, G_3756GAT_OUT, G_3755GAT_OUT, G_3751GAT_OUT, 
      G_3748GAT_OUT, G_3747GAT_OUT, G_3746GAT_OUT, G_3742GAT_OUT, G_3739GAT_OUT
      , G_3736GAT_OUT, G_3735GAT_OUT, G_3734GAT_OUT, G_3730GAT_OUT, 
      G_3727GAT_OUT, G_3724GAT_OUT, G_3721GAT_OUT, G_3718GAT_OUT, G_3715GAT_OUT
      , G_3712GAT_OUT, G_3709GAT_OUT, G_3706GAT_OUT, G_3702GAT_OUT, 
      G_3699GAT_OUT, G_3698GAT_OUT, G_3697GAT_OUT, G_3693GAT_OUT, G_3690GAT_OUT
      , G_3687GAT_OUT, G_3686GAT_OUT, G_3685GAT_OUT, G_3681GAT_OUT, 
      G_3678GAT_OUT, G_3677GAT_OUT, G_3676GAT_OUT, G_3675GAT_OUT, G_3674GAT_OUT
      , G_3673GAT_OUT, G_3672GAT_OUT, G_3671GAT_OUT, G_3670GAT_OUT, 
      G_3669GAT_OUT, G_3668GAT_OUT, G_3667GAT_OUT, G_3666GAT_OUT, G_3665GAT_OUT
      , G_3664GAT_OUT, G_3663GAT_OUT, G_3662GAT_OUT, G_3659GAT_OUT, 
      G_3658GAT_OUT, G_3657GAT_OUT, G_3653GAT_OUT, G_3650GAT_OUT, G_3647GAT_OUT
      , G_3646GAT_OUT, G_3645GAT_OUT, G_3641GAT_OUT, G_3638GAT_OUT, 
      G_3637GAT_OUT, G_3636GAT_OUT, G_3632GAT_OUT, G_3628GAT_OUT, G_3624GAT_OUT
      , G_3620GAT_OUT, G_3616GAT_OUT, G_3612GAT_OUT, G_3608GAT_OUT, 
      G_3604GAT_OUT, G_3603GAT_OUT, G_3602GAT_OUT, G_3598GAT_OUT, G_3595GAT_OUT
      , G_3592GAT_OUT, G_3591GAT_OUT, G_3590GAT_OUT, G_3586GAT_OUT, 
      G_3583GAT_OUT, G_3582GAT_OUT, G_3581GAT_OUT, G_3577GAT_OUT, G_3574GAT_OUT
      , G_3571GAT_OUT, G_3568GAT_OUT, G_3565GAT_OUT, G_3562GAT_OUT, 
      G_3559GAT_OUT, G_3556GAT_OUT, G_3553GAT_OUT, G_3548GAT_OUT, G_3545GAT_OUT
      , G_3542GAT_OUT, G_3541GAT_OUT, G_3540GAT_OUT, G_3536GAT_OUT, 
      G_3533GAT_OUT, G_3532GAT_OUT, G_3531GAT_OUT, G_3527GAT_OUT, G_3524GAT_OUT
      , G_3521GAT_OUT, G_3520GAT_OUT, G_3519GAT_OUT, G_3516GAT_OUT, 
      G_3515GAT_OUT, G_3514GAT_OUT, G_3511GAT_OUT, G_3510GAT_OUT, G_3509GAT_OUT
      , G_3506GAT_OUT, G_3505GAT_OUT, G_3504GAT_OUT, G_3501GAT_OUT, 
      G_3500GAT_OUT, G_3499GAT_OUT, G_3496GAT_OUT, G_3495GAT_OUT, G_3494GAT_OUT
      , G_3491GAT_OUT, G_3490GAT_OUT, G_3489GAT_OUT, G_3486GAT_OUT, 
      G_3485GAT_OUT, G_3484GAT_OUT, G_3481GAT_OUT, G_3480GAT_OUT, G_3479GAT_OUT
      , G_3476GAT_OUT, G_3475GAT_OUT, G_3474GAT_OUT, G_3470GAT_OUT, 
      G_3467GAT_OUT, G_3466GAT_OUT, G_3465GAT_OUT, G_3461GAT_OUT, G_3458GAT_OUT
      , G_3455GAT_OUT, G_3454GAT_OUT, G_3453GAT_OUT, G_3449GAT_OUT, 
      G_3445GAT_OUT, G_3441GAT_OUT, G_3437GAT_OUT, G_3433GAT_OUT, G_3429GAT_OUT
      , G_3425GAT_OUT, G_3421GAT_OUT, G_3417GAT_OUT, G_3413GAT_OUT, 
      G_3410GAT_OUT, G_3409GAT_OUT, G_3408GAT_OUT, G_3404GAT_OUT, G_3401GAT_OUT
      , G_3398GAT_OUT, G_3397GAT_OUT, G_3396GAT_OUT, G_3392GAT_OUT, 
      G_3389GAT_OUT, G_3386GAT_OUT, G_3383GAT_OUT, G_3380GAT_OUT, G_3377GAT_OUT
      , G_3374GAT_OUT, G_3371GAT_OUT, G_3368GAT_OUT, G_3365GAT_OUT, 
      G_3362GAT_OUT, G_3361GAT_OUT, G_3360GAT_OUT, G_3356GAT_OUT, G_3353GAT_OUT
      , G_3350GAT_OUT, G_3349GAT_OUT, G_3348GAT_OUT, G_3344GAT_OUT, 
      G_3341GAT_OUT, G_3340GAT_OUT, G_3339GAT_OUT, G_3338GAT_OUT, G_3337GAT_OUT
      , G_3336GAT_OUT, G_3335GAT_OUT, G_3334GAT_OUT, G_3333GAT_OUT, 
      G_3332GAT_OUT, G_3331GAT_OUT, G_3330GAT_OUT, G_3329GAT_OUT, G_3328GAT_OUT
      , G_3327GAT_OUT, G_3326GAT_OUT, G_3325GAT_OUT, G_3324GAT_OUT, 
      G_3323GAT_OUT, G_3322GAT_OUT, G_3321GAT_OUT, G_3317GAT_OUT, G_3314GAT_OUT
      , G_3311GAT_OUT, G_3310GAT_OUT, G_3309GAT_OUT, G_3305GAT_OUT, 
      G_3302GAT_OUT, G_3301GAT_OUT, G_3300GAT_OUT, G_3296GAT_OUT, G_3292GAT_OUT
      , G_3288GAT_OUT, G_3284GAT_OUT, G_3280GAT_OUT, G_3276GAT_OUT, 
      G_3272GAT_OUT, G_3268GAT_OUT, G_3264GAT_OUT, G_3260GAT_OUT, G_3257GAT_OUT
      , G_3254GAT_OUT, G_3253GAT_OUT, G_3252GAT_OUT, G_3248GAT_OUT, 
      G_3245GAT_OUT, G_3244GAT_OUT, G_3243GAT_OUT, G_3239GAT_OUT, G_3236GAT_OUT
      , G_3233GAT_OUT, G_3230GAT_OUT, G_3227GAT_OUT, G_3224GAT_OUT, 
      G_3221GAT_OUT, G_3218GAT_OUT, G_3215GAT_OUT, G_3212GAT_OUT, G_3208GAT_OUT
      , G_3207GAT_OUT, G_3206GAT_OUT, G_3202GAT_OUT, G_3199GAT_OUT, 
      G_3198GAT_OUT, G_3197GAT_OUT, G_3193GAT_OUT, G_3190GAT_OUT, G_3187GAT_OUT
      , G_3186GAT_OUT, G_3185GAT_OUT, G_3182GAT_OUT, G_3181GAT_OUT, 
      G_3180GAT_OUT, G_3177GAT_OUT, G_3176GAT_OUT, G_3175GAT_OUT, G_3172GAT_OUT
      , G_3171GAT_OUT, G_3170GAT_OUT, G_3167GAT_OUT, G_3166GAT_OUT, 
      G_3165GAT_OUT, G_3162GAT_OUT, G_3161GAT_OUT, G_3160GAT_OUT, G_3157GAT_OUT
      , G_3156GAT_OUT, G_3155GAT_OUT, G_3152GAT_OUT, G_3151GAT_OUT, 
      G_3150GAT_OUT, G_3147GAT_OUT, G_3146GAT_OUT, G_3145GAT_OUT, G_3142GAT_OUT
      , G_3141GAT_OUT, G_3140GAT_OUT, G_3136GAT_OUT, G_3133GAT_OUT, 
      G_3132GAT_OUT, G_3131GAT_OUT, G_3127GAT_OUT, G_3124GAT_OUT, G_3121GAT_OUT
      , G_3120GAT_OUT, G_3119GAT_OUT, G_3115GAT_OUT, G_3111GAT_OUT, 
      G_3107GAT_OUT, G_3103GAT_OUT, G_3099GAT_OUT, G_3095GAT_OUT, G_3091GAT_OUT
      , G_3087GAT_OUT, G_3083GAT_OUT, G_3079GAT_OUT, G_3076GAT_OUT, 
      G_3075GAT_OUT, G_3074GAT_OUT, G_3070GAT_OUT, G_3067GAT_OUT, G_3064GAT_OUT
      , G_3063GAT_OUT, G_3062GAT_OUT, G_3058GAT_OUT, G_3055GAT_OUT, 
      G_3052GAT_OUT, G_3049GAT_OUT, G_3046GAT_OUT, G_3043GAT_OUT, G_3040GAT_OUT
      , G_3037GAT_OUT, G_3034GAT_OUT, G_3031GAT_OUT, G_3028GAT_OUT, 
      G_3027GAT_OUT, G_3026GAT_OUT, G_3022GAT_OUT, G_3019GAT_OUT, G_3016GAT_OUT
      , G_3015GAT_OUT, G_3014GAT_OUT, G_3010GAT_OUT, G_3007GAT_OUT, 
      G_3006GAT_OUT, G_3005GAT_OUT, G_3004GAT_OUT, G_3003GAT_OUT, G_3002GAT_OUT
      , G_3001GAT_OUT, G_3000GAT_OUT, G_2999GAT_OUT, G_2998GAT_OUT, 
      G_2997GAT_OUT, G_2996GAT_OUT, G_2995GAT_OUT, G_2994GAT_OUT, G_2993GAT_OUT
      , G_2992GAT_OUT, G_2991GAT_OUT, G_2990GAT_OUT, G_2989GAT_OUT, 
      G_2988GAT_OUT, G_2987GAT_OUT, G_2983GAT_OUT, G_2980GAT_OUT, G_2977GAT_OUT
      , G_2976GAT_OUT, G_2975GAT_OUT, G_2971GAT_OUT, G_2968GAT_OUT, 
      G_2967GAT_OUT, G_2966GAT_OUT, G_2962GAT_OUT, G_2958GAT_OUT, G_2954GAT_OUT
      , G_2950GAT_OUT, G_2946GAT_OUT, G_2942GAT_OUT, G_2938GAT_OUT, 
      G_2934GAT_OUT, G_2930GAT_OUT, G_2926GAT_OUT, G_2923GAT_OUT, G_2922GAT_OUT
      , G_2921GAT_OUT, G_2917GAT_OUT, G_2914GAT_OUT, G_2913GAT_OUT, 
      G_2912GAT_OUT, G_2908GAT_OUT, G_2905GAT_OUT, G_2902GAT_OUT, G_2899GAT_OUT
      , G_2896GAT_OUT, G_2893GAT_OUT, G_2890GAT_OUT, G_2887GAT_OUT, 
      G_2884GAT_OUT, G_2881GAT_OUT, G_2878GAT_OUT, G_2873GAT_OUT, G_2870GAT_OUT
      , G_2869GAT_OUT, G_2868GAT_OUT, G_2864GAT_OUT, G_2861GAT_OUT, 
      G_2858GAT_OUT, G_2857GAT_OUT, G_2856GAT_OUT, G_2853GAT_OUT, G_2852GAT_OUT
      , G_2851GAT_OUT, G_2848GAT_OUT, G_2847GAT_OUT, G_2846GAT_OUT, 
      G_2843GAT_OUT, G_2842GAT_OUT, G_2841GAT_OUT, G_2838GAT_OUT, G_2837GAT_OUT
      , G_2836GAT_OUT, G_2833GAT_OUT, G_2832GAT_OUT, G_2831GAT_OUT, 
      G_2828GAT_OUT, G_2827GAT_OUT, G_2826GAT_OUT, G_2823GAT_OUT, G_2822GAT_OUT
      , G_2821GAT_OUT, G_2818GAT_OUT, G_2817GAT_OUT, G_2816GAT_OUT, 
      G_2813GAT_OUT, G_2812GAT_OUT, G_2811GAT_OUT, G_2808GAT_OUT, G_2807GAT_OUT
      , G_2806GAT_OUT, G_2803GAT_OUT, G_2802GAT_OUT, G_2801GAT_OUT, 
      G_2797GAT_OUT, G_2794GAT_OUT, G_2791GAT_OUT, G_2790GAT_OUT, G_2789GAT_OUT
      , G_2785GAT_OUT, G_2781GAT_OUT, G_2777GAT_OUT, G_2773GAT_OUT, 
      G_2769GAT_OUT, G_2765GAT_OUT, G_2761GAT_OUT, G_2757GAT_OUT, G_2753GAT_OUT
      , G_2749GAT_OUT, G_2745GAT_OUT, G_2744GAT_OUT, G_2743GAT_OUT, 
      G_2739GAT_OUT, G_2736GAT_OUT, G_2733GAT_OUT, G_2732GAT_OUT, G_2731GAT_OUT
      , G_2727GAT_OUT, G_2724GAT_OUT, G_2721GAT_OUT, G_2718GAT_OUT, 
      G_2715GAT_OUT, G_2712GAT_OUT, G_2709GAT_OUT, G_2706GAT_OUT, G_2703GAT_OUT
      , G_2700GAT_OUT, G_2697GAT_OUT, G_2694GAT_OUT, G_2690GAT_OUT, 
      G_2687GAT_OUT, G_2684GAT_OUT, G_2683GAT_OUT, G_2682GAT_OUT, G_2678GAT_OUT
      , G_2675GAT_OUT, G_2674GAT_OUT, G_2673GAT_OUT, G_2672GAT_OUT, 
      G_2671GAT_OUT, G_2670GAT_OUT, G_2669GAT_OUT, G_2668GAT_OUT, G_2667GAT_OUT
      , G_2666GAT_OUT, G_2665GAT_OUT, G_2664GAT_OUT, G_2663GAT_OUT, 
      G_2662GAT_OUT, G_2661GAT_OUT, G_2660GAT_OUT, G_2659GAT_OUT, G_2658GAT_OUT
      , G_2657GAT_OUT, G_2656GAT_OUT, G_2655GAT_OUT, G_2654GAT_OUT, 
      G_2653GAT_OUT, G_2650GAT_OUT, G_2649GAT_OUT, G_2648GAT_OUT, G_2644GAT_OUT
      , G_2641GAT_OUT, G_2640GAT_OUT, G_2639GAT_OUT, G_2635GAT_OUT, 
      G_2631GAT_OUT, G_2627GAT_OUT, G_2623GAT_OUT, G_2619GAT_OUT, G_2615GAT_OUT
      , G_2611GAT_OUT, G_2607GAT_OUT, G_2603GAT_OUT, G_2599GAT_OUT, 
      G_2595GAT_OUT, G_2591GAT_OUT, G_2588GAT_OUT, G_2587GAT_OUT, G_2586GAT_OUT
      , G_2582GAT_OUT, G_2579GAT_OUT, G_2576GAT_OUT, G_2573GAT_OUT, 
      G_2570GAT_OUT, G_2567GAT_OUT, G_2564GAT_OUT, G_2561GAT_OUT, G_2558GAT_OUT
      , G_2555GAT_OUT, G_2552GAT_OUT, G_2549GAT_OUT, G_2545GAT_OUT, 
      G_2544GAT_OUT, G_2543GAT_OUT, G_2539GAT_OUT, G_2536GAT_OUT, G_2533GAT_OUT
      , G_2532GAT_OUT, G_2531GAT_OUT, G_2528GAT_OUT, G_2527GAT_OUT, 
      G_2526GAT_OUT, G_2523GAT_OUT, G_2522GAT_OUT, G_2521GAT_OUT, G_2518GAT_OUT
      , G_2517GAT_OUT, G_2516GAT_OUT, G_2513GAT_OUT, G_2512GAT_OUT, 
      G_2511GAT_OUT, G_2508GAT_OUT, G_2507GAT_OUT, G_2506GAT_OUT, G_2503GAT_OUT
      , G_2502GAT_OUT, G_2501GAT_OUT, G_2498GAT_OUT, G_2497GAT_OUT, 
      G_2496GAT_OUT, G_2493GAT_OUT, G_2492GAT_OUT, G_2491GAT_OUT, G_2488GAT_OUT
      , G_2487GAT_OUT, G_2486GAT_OUT, G_2483GAT_OUT, G_2482GAT_OUT, 
      G_2481GAT_OUT, G_2478GAT_OUT, G_2477GAT_OUT, G_2476GAT_OUT, G_2475GAT_OUT
      , G_2474GAT_OUT, G_2470GAT_OUT, G_2467GAT_OUT, G_2464GAT_OUT, 
      G_2463GAT_OUT, G_2462GAT_OUT, G_2458GAT_OUT, G_2454GAT_OUT, G_2450GAT_OUT
      , G_2446GAT_OUT, G_2442GAT_OUT, G_2438GAT_OUT, G_2434GAT_OUT, 
      G_2430GAT_OUT, G_2426GAT_OUT, G_2422GAT_OUT, G_2418GAT_OUT, G_2414GAT_OUT
      , G_2410GAT_OUT, G_2407GAT_OUT, G_2404GAT_OUT, G_2403GAT_OUT, 
      G_2402GAT_OUT, G_2398GAT_OUT, G_2395GAT_OUT, G_2392GAT_OUT, G_2389GAT_OUT
      , G_2386GAT_OUT, G_2383GAT_OUT, G_2380GAT_OUT, G_2377GAT_OUT, 
      G_2374GAT_OUT, G_2371GAT_OUT, G_2368GAT_OUT, G_2365GAT_OUT, G_2362GAT_OUT
      , G_2359GAT_OUT, G_2358GAT_OUT, G_2357GAT_OUT, G_2353GAT_OUT, 
      G_2350GAT_OUT, G_2349GAT_OUT, G_2348GAT_OUT, G_2347GAT_OUT, G_2346GAT_OUT
      , G_2345GAT_OUT, G_2344GAT_OUT, G_2343GAT_OUT, G_2342GAT_OUT, 
      G_2341GAT_OUT, G_2340GAT_OUT, G_2339GAT_OUT, G_2338GAT_OUT, G_2337GAT_OUT
      , G_2336GAT_OUT, G_2335GAT_OUT, G_2334GAT_OUT, G_2333GAT_OUT, 
      G_2332GAT_OUT, G_2331GAT_OUT, G_2330GAT_OUT, G_2329GAT_OUT, G_2328GAT_OUT
      , G_2327GAT_OUT, G_2326GAT_OUT, G_2322GAT_OUT, G_2319GAT_OUT, 
      G_2318GAT_OUT, G_2317GAT_OUT, G_2313GAT_OUT, G_2309GAT_OUT, G_2305GAT_OUT
      , G_2301GAT_OUT, G_2297GAT_OUT, G_2293GAT_OUT, G_2289GAT_OUT, 
      G_2285GAT_OUT, G_2281GAT_OUT, G_2277GAT_OUT, G_2273GAT_OUT, G_2269GAT_OUT
      , G_2266GAT_OUT, G_2265GAT_OUT, G_2264GAT_OUT, G_2260GAT_OUT, 
      G_2257GAT_OUT, G_2254GAT_OUT, G_2251GAT_OUT, G_2248GAT_OUT, G_2245GAT_OUT
      , G_2242GAT_OUT, G_2239GAT_OUT, G_2236GAT_OUT, G_2233GAT_OUT, 
      G_2230GAT_OUT, G_2227GAT_OUT, G_2224GAT_OUT, G_2222GAT_OUT, G_2221GAT_OUT
      , G_2217GAT_OUT, G_2214GAT_OUT, G_2211GAT_OUT, G_2210GAT_OUT, 
      G_2209GAT_OUT, G_2206GAT_OUT, G_2205GAT_OUT, G_2204GAT_OUT, G_2201GAT_OUT
      , G_2200GAT_OUT, G_2199GAT_OUT, G_2196GAT_OUT, G_2195GAT_OUT, 
      G_2194GAT_OUT, G_2191GAT_OUT, G_2190GAT_OUT, G_2189GAT_OUT, G_2186GAT_OUT
      , G_2185GAT_OUT, G_2184GAT_OUT, G_2181GAT_OUT, G_2180GAT_OUT, 
      G_2179GAT_OUT, G_2176GAT_OUT, G_2175GAT_OUT, G_2174GAT_OUT, G_2171GAT_OUT
      , G_2170GAT_OUT, G_2169GAT_OUT, G_2166GAT_OUT, G_2165GAT_OUT, 
      G_2164GAT_OUT, G_2161GAT_OUT, G_2160GAT_OUT, G_2159GAT_OUT, G_2156GAT_OUT
      , G_2155GAT_OUT, G_2154GAT_OUT, G_2151GAT_OUT, G_2150GAT_OUT, 
      G_2149GAT_OUT, G_2145GAT_OUT, G_2142GAT_OUT, G_2139GAT_OUT, G_2138GAT_OUT
      , G_2137GAT_OUT, G_2133GAT_OUT, G_2129GAT_OUT, G_2125GAT_OUT, 
      G_2121GAT_OUT, G_2117GAT_OUT, G_2113GAT_OUT, G_2109GAT_OUT, G_2105GAT_OUT
      , G_2101GAT_OUT, G_2097GAT_OUT, G_2093GAT_OUT, G_2089GAT_OUT, 
      G_2085GAT_OUT, G_2082GAT_OUT, G_2081GAT_OUT, G_2080GAT_OUT, G_2076GAT_OUT
      , G_2073GAT_OUT, G_2070GAT_OUT, G_2067GAT_OUT, G_2064GAT_OUT, 
      G_2061GAT_OUT, G_2058GAT_OUT, G_2055GAT_OUT, G_2052GAT_OUT, G_2049GAT_OUT
      , G_2046GAT_OUT, G_2043GAT_OUT, G_2040GAT_OUT, G_2037GAT_OUT, 
      G_2033GAT_OUT, G_2030GAT_OUT, G_2029GAT_OUT, G_2028GAT_OUT, G_2027GAT_OUT
      , G_2026GAT_OUT, G_2025GAT_OUT, G_2024GAT_OUT, G_2023GAT_OUT, 
      G_2022GAT_OUT, G_2021GAT_OUT, G_2020GAT_OUT, G_2019GAT_OUT, G_2018GAT_OUT
      , G_2017GAT_OUT, G_2016GAT_OUT, G_2015GAT_OUT, G_2014GAT_OUT, 
      G_2013GAT_OUT, G_2012GAT_OUT, G_2011GAT_OUT, G_2010GAT_OUT, G_2009GAT_OUT
      , G_2008GAT_OUT, G_2007GAT_OUT, G_2006GAT_OUT, G_2005GAT_OUT, 
      G_2004GAT_OUT, G_2001GAT_OUT, G_2000GAT_OUT, G_1999GAT_OUT, G_1995GAT_OUT
      , G_1991GAT_OUT, G_1987GAT_OUT, G_1983GAT_OUT, G_1979GAT_OUT, 
      G_1975GAT_OUT, G_1971GAT_OUT, G_1967GAT_OUT, G_1963GAT_OUT, G_1959GAT_OUT
      , G_1955GAT_OUT, G_1951GAT_OUT, G_1947GAT_OUT, G_1946GAT_OUT, 
      G_1945GAT_OUT, G_1941GAT_OUT, G_1938GAT_OUT, G_1935GAT_OUT, G_1932GAT_OUT
      , G_1929GAT_OUT, G_1926GAT_OUT, G_1923GAT_OUT, G_1920GAT_OUT, 
      G_1917GAT_OUT, G_1914GAT_OUT, G_1911GAT_OUT, G_1908GAT_OUT, G_1905GAT_OUT
      , G_1902GAT_OUT, G_1897GAT_OUT, G_1894GAT_OUT, G_1891GAT_OUT, 
      G_1890GAT_OUT, G_1889GAT_OUT, G_1886GAT_OUT, G_1885GAT_OUT, G_1884GAT_OUT
      , G_1881GAT_OUT, G_1880GAT_OUT, G_1879GAT_OUT, G_1876GAT_OUT, 
      G_1875GAT_OUT, G_1874GAT_OUT, G_1871GAT_OUT, G_1870GAT_OUT, G_1869GAT_OUT
      , G_1866GAT_OUT, G_1865GAT_OUT, G_1864GAT_OUT, G_1861GAT_OUT, 
      G_1860GAT_OUT, G_1859GAT_OUT, G_1856GAT_OUT, G_1855GAT_OUT, G_1854GAT_OUT
      , G_1851GAT_OUT, G_1850GAT_OUT, G_1849GAT_OUT, G_1846GAT_OUT, 
      G_1845GAT_OUT, G_1844GAT_OUT, G_1841GAT_OUT, G_1840GAT_OUT, G_1839GAT_OUT
      , G_1836GAT_OUT, G_1835GAT_OUT, G_1834GAT_OUT, G_1831GAT_OUT, 
      G_1830GAT_OUT, G_1829GAT_OUT, G_1826GAT_OUT, G_1825GAT_OUT, G_1824GAT_OUT
      , G_1821GAT_OUT, G_1820GAT_OUT, G_1819GAT_OUT, G_1815GAT_OUT, 
      G_1811GAT_OUT, G_1807GAT_OUT, G_1803GAT_OUT, G_1799GAT_OUT, G_1795GAT_OUT
      , G_1791GAT_OUT, G_1787GAT_OUT, G_1783GAT_OUT, G_1779GAT_OUT, 
      G_1775GAT_OUT, G_1771GAT_OUT, G_1767GAT_OUT, G_1763GAT_OUT, G_1759GAT_OUT
      , G_1756GAT_OUT, G_1753GAT_OUT, G_1750GAT_OUT, G_1747GAT_OUT, 
      G_1744GAT_OUT, G_1741GAT_OUT, G_1738GAT_OUT, G_1735GAT_OUT, G_1732GAT_OUT
      , G_1729GAT_OUT, G_1726GAT_OUT, G_1723GAT_OUT, G_1720GAT_OUT, 
      G_1717GAT_OUT, G_1714GAT_OUT, G_1713GAT_OUT, G_1712GAT_OUT, G_1711GAT_OUT
      , G_1710GAT_OUT, G_1709GAT_OUT, G_1708GAT_OUT, G_1707GAT_OUT, 
      G_1706GAT_OUT, G_1705GAT_OUT, G_1704GAT_OUT, G_1703GAT_OUT, G_1702GAT_OUT
      , G_1701GAT_OUT, G_1700GAT_OUT, G_1699GAT_OUT, G_1698GAT_OUT, 
      G_1697GAT_OUT, G_1696GAT_OUT, G_1695GAT_OUT, G_1694GAT_OUT, G_1693GAT_OUT
      , G_1692GAT_OUT, G_1691GAT_OUT, G_1690GAT_OUT, G_1689GAT_OUT, 
      G_1688GAT_OUT, G_1687GAT_OUT, G_1686GAT_OUT, G_1685GAT_OUT, G_1684GAT_OUT
      , G_1680GAT_OUT, G_1676GAT_OUT, G_1672GAT_OUT, G_1668GAT_OUT, 
      G_1664GAT_OUT, G_1660GAT_OUT, G_1656GAT_OUT, G_1652GAT_OUT, G_1648GAT_OUT
      , G_1644GAT_OUT, G_1640GAT_OUT, G_1636GAT_OUT, G_1632GAT_OUT, 
      G_1628GAT_OUT, G_1624GAT_OUT, G_1621GAT_OUT, G_1618GAT_OUT, G_1615GAT_OUT
      , G_1612GAT_OUT, G_1609GAT_OUT, G_1606GAT_OUT, G_1603GAT_OUT, 
      G_1600GAT_OUT, G_1597GAT_OUT, G_1594GAT_OUT, G_1591GAT_OUT, G_1588GAT_OUT
      , G_1585GAT_OUT, G_1582GAT_OUT, G_1578GAT_OUT, G_1577GAT_OUT, 
      G_1576GAT_OUT, G_1573GAT_OUT, G_1572GAT_OUT, G_1571GAT_OUT, G_1568GAT_OUT
      , G_1567GAT_OUT, G_1566GAT_OUT, G_1563GAT_OUT, G_1562GAT_OUT, 
      G_1561GAT_OUT, G_1558GAT_OUT, G_1557GAT_OUT, G_1556GAT_OUT, G_1553GAT_OUT
      , G_1552GAT_OUT, G_1551GAT_OUT, G_1548GAT_OUT, G_1547GAT_OUT, 
      G_1546GAT_OUT, G_1543GAT_OUT, G_1542GAT_OUT, G_1541GAT_OUT, G_1538GAT_OUT
      , G_1537GAT_OUT, G_1536GAT_OUT, G_1533GAT_OUT, G_1532GAT_OUT, 
      G_1531GAT_OUT, G_1528GAT_OUT, G_1527GAT_OUT, G_1526GAT_OUT, G_1523GAT_OUT
      , G_1522GAT_OUT, G_1521GAT_OUT, G_1518GAT_OUT, G_1517GAT_OUT, 
      G_1516GAT_OUT, G_1513GAT_OUT, G_1512GAT_OUT, G_1511GAT_OUT, G_1508GAT_OUT
      , G_1507GAT_OUT, G_1506GAT_OUT, G_1502GAT_OUT, G_1498GAT_OUT, 
      G_1494GAT_OUT, G_1490GAT_OUT, G_1486GAT_OUT, G_1482GAT_OUT, G_1478GAT_OUT
      , G_1474GAT_OUT, G_1470GAT_OUT, G_1466GAT_OUT, G_1462GAT_OUT, 
      G_1458GAT_OUT, G_1454GAT_OUT, G_1450GAT_OUT, G_1446GAT_OUT, G_1443GAT_OUT
      , G_1440GAT_OUT, G_1437GAT_OUT, G_1434GAT_OUT, G_1431GAT_OUT, 
      G_1428GAT_OUT, G_1425GAT_OUT, G_1422GAT_OUT, G_1419GAT_OUT, G_1416GAT_OUT
      , G_1413GAT_OUT, G_1410GAT_OUT, G_1407GAT_OUT, G_1404GAT_OUT, 
      G_1401GAT_OUT, G_1400GAT_OUT, G_1399GAT_OUT, G_1398GAT_OUT, G_1397GAT_OUT
      , G_1396GAT_OUT, G_1395GAT_OUT, G_1394GAT_OUT, G_1393GAT_OUT, 
      G_1392GAT_OUT, G_1391GAT_OUT, G_1390GAT_OUT, G_1389GAT_OUT, G_1388GAT_OUT
      , G_1387GAT_OUT, G_1386GAT_OUT, G_1385GAT_OUT, G_1384GAT_OUT, 
      G_1383GAT_OUT, G_1382GAT_OUT, G_1381GAT_OUT, G_1380GAT_OUT, G_1379GAT_OUT
      , G_1378GAT_OUT, G_1377GAT_OUT, G_1376GAT_OUT, G_1375GAT_OUT, 
      G_1374GAT_OUT, G_1373GAT_OUT, G_1372GAT_OUT, G_1371GAT_OUT, G_1367GAT_OUT
      , G_1363GAT_OUT, G_1359GAT_OUT, G_1355GAT_OUT, G_1351GAT_OUT, 
      G_1347GAT_OUT, G_1343GAT_OUT, G_1339GAT_OUT, G_1335GAT_OUT, G_1331GAT_OUT
      , G_1327GAT_OUT, G_1323GAT_OUT, G_1319GAT_OUT, G_1315GAT_OUT, 
      G_1311GAT_OUT, G_1308GAT_OUT, G_1305GAT_OUT, G_1302GAT_OUT, G_1299GAT_OUT
      , G_1296GAT_OUT, G_1293GAT_OUT, G_1290GAT_OUT, G_1287GAT_OUT, 
      G_1284GAT_OUT, G_1281GAT_OUT, G_1278GAT_OUT, G_1275GAT_OUT, G_1272GAT_OUT
      , G_1269GAT_OUT, G_1266GAT_OUT, G_1263GAT_OUT, G_1260GAT_OUT, 
      G_1257GAT_OUT, G_1254GAT_OUT, G_1251GAT_OUT, G_1248GAT_OUT, G_1245GAT_OUT
      , G_1242GAT_OUT, G_1239GAT_OUT, G_1236GAT_OUT, G_1233GAT_OUT, 
      G_1230GAT_OUT, G_1227GAT_OUT, G_1224GAT_OUT, G_1221GAT_OUT, G_1218GAT_OUT
      , G_1215GAT_OUT, G_1212GAT_OUT, G_1209GAT_OUT, G_1206GAT_OUT, 
      G_1203GAT_OUT, G_1200GAT_OUT, G_1197GAT_OUT, G_1194GAT_OUT, G_1191GAT_OUT
      , G_1188GAT_OUT, G_1185GAT_OUT, G_1182GAT_OUT, G_1179GAT_OUT, 
      G_1176GAT_OUT, G_1173GAT_OUT, G_1170GAT_OUT, G_1167GAT_OUT, G_1164GAT_OUT
      , G_1161GAT_OUT, G_1158GAT_OUT, G_1155GAT_OUT, G_1152GAT_OUT, 
      G_1149GAT_OUT, G_1146GAT_OUT, G_1143GAT_OUT, G_1140GAT_OUT, G_1137GAT_OUT
      , G_1134GAT_OUT, G_1131GAT_OUT, G_1128GAT_OUT, G_1125GAT_OUT, 
      G_1122GAT_OUT, G_1119GAT_OUT, G_1116GAT_OUT, G_1113GAT_OUT, G_1110GAT_OUT
      , G_1107GAT_OUT, G_1104GAT_OUT, G_1101GAT_OUT, G_1098GAT_OUT, 
      G_1095GAT_OUT, G_1092GAT_OUT, G_1089GAT_OUT, G_1086GAT_OUT, G_1083GAT_OUT
      , G_1080GAT_OUT, G_1077GAT_OUT, G_1074GAT_OUT, G_1071GAT_OUT, 
      G_1068GAT_OUT, G_1065GAT_OUT, G_1062GAT_OUT, G_1059GAT_OUT, G_1056GAT_OUT
      , G_1053GAT_OUT, G_1050GAT_OUT, G_1047GAT_OUT, G_1044GAT_OUT, 
      G_1041GAT_OUT, G_1038GAT_OUT, G_1035GAT_OUT, G_1032GAT_OUT, G_1029GAT_OUT
      , G_1026GAT_OUT, G_1023GAT_OUT, G_1020GAT_OUT, G_1017GAT_OUT, 
      G_1014GAT_OUT, G_1011GAT_OUT, G_1008GAT_OUT, G_1005GAT_OUT, G_1002GAT_OUT
      , G_999GAT_OUT, G_996GAT_OUT, G_993GAT_OUT, G_990GAT_OUT, G_987GAT_OUT, 
      G_984GAT_OUT, G_981GAT_OUT, G_978GAT_OUT, G_975GAT_OUT, G_972GAT_OUT, 
      G_969GAT_OUT, G_966GAT_OUT, G_963GAT_OUT, G_960GAT_OUT, G_957GAT_OUT, 
      G_954GAT_OUT, G_951GAT_OUT, G_948GAT_OUT, G_945GAT_OUT, G_942GAT_OUT, 
      G_939GAT_OUT, G_936GAT_OUT, G_933GAT_OUT, G_930GAT_OUT, G_927GAT_OUT, 
      G_924GAT_OUT, G_921GAT_OUT, G_918GAT_OUT, G_915GAT_OUT, G_912GAT_OUT, 
      G_909GAT_OUT, G_906GAT_OUT, G_903GAT_OUT, G_900GAT_OUT, G_897GAT_OUT, 
      G_894GAT_OUT, G_891GAT_OUT, G_888GAT_OUT, G_885GAT_OUT, G_882GAT_OUT, 
      G_879GAT_OUT, G_876GAT_OUT, G_873GAT_OUT, G_870GAT_OUT, G_867GAT_OUT, 
      G_864GAT_OUT, G_861GAT_OUT, G_858GAT_OUT, G_855GAT_OUT, G_852GAT_OUT, 
      G_849GAT_OUT, G_846GAT_OUT, G_843GAT_OUT, G_840GAT_OUT, G_837GAT_OUT, 
      G_834GAT_OUT, G_831GAT_OUT, G_828GAT_OUT, G_825GAT_OUT, G_822GAT_OUT, 
      G_819GAT_OUT, G_816GAT_OUT, G_813GAT_OUT, G_810GAT_OUT, G_807GAT_OUT, 
      G_804GAT_OUT, G_801GAT_OUT, G_798GAT_OUT, G_795GAT_OUT, G_792GAT_OUT, 
      G_789GAT_OUT, G_786GAT_OUT, G_783GAT_OUT, G_780GAT_OUT, G_777GAT_OUT, 
      G_774GAT_OUT, G_771GAT_OUT, G_768GAT_OUT, G_765GAT_OUT, G_762GAT_OUT, 
      G_759GAT_OUT, G_756GAT_OUT, G_753GAT_OUT, G_750GAT_OUT, G_747GAT_OUT, 
      G_744GAT_OUT, G_741GAT_OUT, G_738GAT_OUT, G_735GAT_OUT, G_732GAT_OUT, 
      G_729GAT_OUT, G_726GAT_OUT, G_723GAT_OUT, G_720GAT_OUT, G_717GAT_OUT, 
      G_714GAT_OUT, G_711GAT_OUT, G_708GAT_OUT, G_705GAT_OUT, G_702GAT_OUT, 
      G_699GAT_OUT, G_696GAT_OUT, G_693GAT_OUT, G_690GAT_OUT, G_687GAT_OUT, 
      G_684GAT_OUT, G_681GAT_OUT, G_678GAT_OUT, G_675GAT_OUT, G_672GAT_OUT, 
      G_669GAT_OUT, G_666GAT_OUT, G_663GAT_OUT, G_660GAT_OUT, G_657GAT_OUT, 
      G_654GAT_OUT, G_651GAT_OUT, G_648GAT_OUT, G_645GAT_OUT, G_642GAT_OUT, 
      G_639GAT_OUT, G_636GAT_OUT, G_633GAT_OUT, G_630GAT_OUT, G_627GAT_OUT, 
      G_624GAT_OUT, G_621GAT_OUT, G_618GAT_OUT, G_615GAT_OUT, G_612GAT_OUT, 
      G_609GAT_OUT, G_606GAT_OUT, G_603GAT_OUT, G_600GAT_OUT, G_597GAT_OUT, 
      G_594GAT_OUT, G_591GAT_OUT, G_588GAT_OUT, G_585GAT_OUT, G_582GAT_OUT, 
      G_579GAT_OUT, G_576GAT_OUT, G_573GAT_OUT, G_570GAT_OUT, G_567GAT_OUT, 
      G_564GAT_OUT, G_561GAT_OUT, G_558GAT_OUT, G_555GAT_OUT, G_552GAT_OUT, 
      G_549GAT_OUT, G_546GAT_OUT : std_logic;

begin

G_1GAT <= datai(31);
G_18GAT <= datai(30);
G_35GAT <= datai(29);
G_52GAT <= datai(28);
G_69GAT <= datai(27);
G_86GAT <= datai(26);
G_103GAT <= datai(25);
G_120GAT <= datai(24);
G_137GAT <= datai(23);
G_154GAT <= datai(22);
G_171GAT <= datai(21);
G_188GAT <= datai(20);
G_205GAT <= datai(19);
G_222GAT <= datai(18);
G_239GAT <= datai(17);
G_256GAT <= datai(16);
G_273GAT <= datai(15);
G_290GAT <= datai(14);
G_307GAT <= datai(13);
G_324GAT <= datai(12);
G_341GAT <= datai(11);
G_358GAT <= datai(10);
G_375GAT <= datai(9);
G_392GAT <= datai(8);
G_409GAT <= datai(7);
G_426GAT <= datai(6);
G_443GAT <= datai(5);
G_460GAT <= datai(4);
G_477GAT <= datai(3);
G_494GAT <= datai(2);
G_511GAT <= datai(1);
G_528GAT <= datai(0);


datao(31) <= G_545GAT_PO;
datao(30) <= G_1581GAT_PO;
datao(29) <= G_1901GAT_PO;
datao(28) <= G_2223GAT_PO;
datao(27) <= G_2548GAT_PO;
datao(26) <= G_2877GAT_PO;
datao(25) <= G_3211GAT_PO;
datao(24) <= G_3552GAT_PO;
datao(23) <= G_3895GAT_PO;
datao(22) <= G_4241GAT_PO;
datao(21) <= G_4591GAT_PO;
datao(20) <= G_4946GAT_PO;
datao(19) <= G_5308GAT_PO;
datao(18) <= G_5672GAT_PO;
datao(17) <= G_5971GAT_PO;
datao(16) <= G_6123GAT_PO;
datao(15) <= G_6150GAT_PO;
datao(14) <= G_6160GAT_PO;
datao(13) <= G_6170GAT_PO;
datao(12) <= G_6180GAT_PO;
datao(11) <= G_6190GAT_PO;
datao(10) <= G_6200GAT_PO;
datao(9) <= G_6210GAT_PO;
datao(8) <= G_6220GAT_PO;
datao(7) <= G_6230GAT_PO;
datao(6) <= G_6240GAT_PO;
datao(5) <= G_6250GAT_PO;
datao(4) <= G_6260GAT_PO;
datao(3) <= G_6270GAT_PO;
datao(2) <= G_6280GAT_PO;
datao(1) <= G_6287GAT_PO;
datao(0) <= G_6288GAT_PO;







   
   G_6286GAT : Nor_gate port map( I1 => G_6281GAT_OUT, I2 => G_6277GAT_OUT, O 
                           => G_6286GAT_OUT);
   G_6285GAT : Nor_gate port map( I1 => G_5727GAT_OUT, I2 => G_6281GAT_OUT, O 
                           => G_6285GAT_OUT);
   G_6281GAT : Nor_gate port map( I1 => G_5727GAT_OUT, I2 => G_6277GAT_OUT, O 
                           => G_6281GAT_OUT);
   G_6277GAT : Nor_gate port map( I1 => G_5666GAT_OUT, I2 => G_6271GAT_OUT, O 
                           => G_6277GAT_OUT);
   G_6276GAT : Nor_gate port map( I1 => G_6271GAT_OUT, I2 => G_6267GAT_OUT, O 
                           => G_6276GAT_OUT);
   G_6275GAT : Nor_gate port map( I1 => G_5782GAT_OUT, I2 => G_6271GAT_OUT, O 
                           => G_6275GAT_OUT);
   G_6271GAT : Nor_gate port map( I1 => G_5782GAT_OUT, I2 => G_6267GAT_OUT, O 
                           => G_6271GAT_OUT);
   G_6267GAT : Nor_gate port map( I1 => G_5721GAT_OUT, I2 => G_6261GAT_OUT, O 
                           => G_6267GAT_OUT);
   G_6266GAT : Nor_gate port map( I1 => G_6261GAT_OUT, I2 => G_6257GAT_OUT, O 
                           => G_6266GAT_OUT);
   G_6265GAT : Nor_gate port map( I1 => G_5831GAT_OUT, I2 => G_6261GAT_OUT, O 
                           => G_6265GAT_OUT);
   G_6261GAT : Nor_gate port map( I1 => G_5831GAT_OUT, I2 => G_6257GAT_OUT, O 
                           => G_6261GAT_OUT);
   G_6257GAT : Nor_gate port map( I1 => G_5776GAT_OUT, I2 => G_6251GAT_OUT, O 
                           => G_6257GAT_OUT);
   G_6256GAT : Nor_gate port map( I1 => G_6251GAT_OUT, I2 => G_6247GAT_OUT, O 
                           => G_6256GAT_OUT);
   G_6255GAT : Nor_gate port map( I1 => G_5879GAT_OUT, I2 => G_6251GAT_OUT, O 
                           => G_6255GAT_OUT);
   G_6251GAT : Nor_gate port map( I1 => G_5879GAT_OUT, I2 => G_6247GAT_OUT, O 
                           => G_6251GAT_OUT);
   G_6247GAT : Nor_gate port map( I1 => G_5825GAT_OUT, I2 => G_6241GAT_OUT, O 
                           => G_6247GAT_OUT);
   G_6246GAT : Nor_gate port map( I1 => G_6241GAT_OUT, I2 => G_6237GAT_OUT, O 
                           => G_6246GAT_OUT);
   G_6245GAT : Nor_gate port map( I1 => G_5925GAT_OUT, I2 => G_6241GAT_OUT, O 
                           => G_6245GAT_OUT);
   G_6241GAT : Nor_gate port map( I1 => G_5925GAT_OUT, I2 => G_6237GAT_OUT, O 
                           => G_6241GAT_OUT);
   G_6237GAT : Nor_gate port map( I1 => G_5873GAT_OUT, I2 => G_6231GAT_OUT, O 
                           => G_6237GAT_OUT);
   G_6236GAT : Nor_gate port map( I1 => G_6231GAT_OUT, I2 => G_6227GAT_OUT, O 
                           => G_6236GAT_OUT);
   G_6235GAT : Nor_gate port map( I1 => G_5968GAT_OUT, I2 => G_6231GAT_OUT, O 
                           => G_6235GAT_OUT);
   G_6231GAT : Nor_gate port map( I1 => G_5968GAT_OUT, I2 => G_6227GAT_OUT, O 
                           => G_6231GAT_OUT);
   G_6227GAT : Nor_gate port map( I1 => G_5919GAT_OUT, I2 => G_6221GAT_OUT, O 
                           => G_6227GAT_OUT);
   G_6226GAT : Nor_gate port map( I1 => G_6221GAT_OUT, I2 => G_6217GAT_OUT, O 
                           => G_6226GAT_OUT);
   G_6225GAT : Nor_gate port map( I1 => G_6002GAT_OUT, I2 => G_6221GAT_OUT, O 
                           => G_6225GAT_OUT);
   G_6221GAT : Nor_gate port map( I1 => G_6002GAT_OUT, I2 => G_6217GAT_OUT, O 
                           => G_6221GAT_OUT);
   G_6217GAT : Nor_gate port map( I1 => G_5962GAT_OUT, I2 => G_6211GAT_OUT, O 
                           => G_6217GAT_OUT);
   G_6216GAT : Nor_gate port map( I1 => G_6211GAT_OUT, I2 => G_6207GAT_OUT, O 
                           => G_6216GAT_OUT);
   G_6215GAT : Nor_gate port map( I1 => G_6032GAT_OUT, I2 => G_6211GAT_OUT, O 
                           => G_6215GAT_OUT);
   G_6211GAT : Nor_gate port map( I1 => G_6032GAT_OUT, I2 => G_6207GAT_OUT, O 
                           => G_6211GAT_OUT);
   G_6207GAT : Nor_gate port map( I1 => G_5996GAT_OUT, I2 => G_6201GAT_OUT, O 
                           => G_6207GAT_OUT);
   G_6206GAT : Nor_gate port map( I1 => G_6201GAT_OUT, I2 => G_6197GAT_OUT, O 
                           => G_6206GAT_OUT);
   G_6205GAT : Nor_gate port map( I1 => G_6058GAT_OUT, I2 => G_6201GAT_OUT, O 
                           => G_6205GAT_OUT);
   G_6201GAT : Nor_gate port map( I1 => G_6058GAT_OUT, I2 => G_6197GAT_OUT, O 
                           => G_6201GAT_OUT);
   G_6197GAT : Nor_gate port map( I1 => G_6026GAT_OUT, I2 => G_6191GAT_OUT, O 
                           => G_6197GAT_OUT);
   G_6196GAT : Nor_gate port map( I1 => G_6191GAT_OUT, I2 => G_6187GAT_OUT, O 
                           => G_6196GAT_OUT);
   G_6195GAT : Nor_gate port map( I1 => G_6082GAT_OUT, I2 => G_6191GAT_OUT, O 
                           => G_6195GAT_OUT);
   G_6191GAT : Nor_gate port map( I1 => G_6082GAT_OUT, I2 => G_6187GAT_OUT, O 
                           => G_6191GAT_OUT);
   G_6187GAT : Nor_gate port map( I1 => G_6052GAT_OUT, I2 => G_6181GAT_OUT, O 
                           => G_6187GAT_OUT);
   G_6186GAT : Nor_gate port map( I1 => G_6181GAT_OUT, I2 => G_6177GAT_OUT, O 
                           => G_6186GAT_OUT);
   G_6185GAT : Nor_gate port map( I1 => G_6103GAT_OUT, I2 => G_6181GAT_OUT, O 
                           => G_6185GAT_OUT);
   G_6181GAT : Nor_gate port map( I1 => G_6103GAT_OUT, I2 => G_6177GAT_OUT, O 
                           => G_6181GAT_OUT);
   G_6177GAT : Nor_gate port map( I1 => G_6076GAT_OUT, I2 => G_6171GAT_OUT, O 
                           => G_6177GAT_OUT);
   G_6176GAT : Nor_gate port map( I1 => G_6171GAT_OUT, I2 => G_6167GAT_OUT, O 
                           => G_6176GAT_OUT);
   G_6175GAT : Nor_gate port map( I1 => G_6120GAT_OUT, I2 => G_6171GAT_OUT, O 
                           => G_6175GAT_OUT);
   G_6171GAT : Nor_gate port map( I1 => G_6120GAT_OUT, I2 => G_6167GAT_OUT, O 
                           => G_6171GAT_OUT);
   G_6167GAT : Nor_gate port map( I1 => G_6097GAT_OUT, I2 => G_6161GAT_OUT, O 
                           => G_6167GAT_OUT);
   G_6166GAT : Nor_gate port map( I1 => G_6161GAT_OUT, I2 => G_6157GAT_OUT, O 
                           => G_6166GAT_OUT);
   G_6165GAT : Nor_gate port map( I1 => G_6130GAT_OUT, I2 => G_6161GAT_OUT, O 
                           => G_6165GAT_OUT);
   G_6161GAT : Nor_gate port map( I1 => G_6130GAT_OUT, I2 => G_6157GAT_OUT, O 
                           => G_6161GAT_OUT);
   G_6157GAT : Nor_gate port map( I1 => G_6114GAT_OUT, I2 => G_6151GAT_OUT, O 
                           => G_6157GAT_OUT);
   G_6156GAT : Nor_gate port map( I1 => G_6151GAT_OUT, I2 => G_6147GAT_OUT, O 
                           => G_6156GAT_OUT);
   G_6155GAT : Nor_gate port map( I1 => G_6135GAT_OUT, I2 => G_6151GAT_OUT, O 
                           => G_6155GAT_OUT);
   G_6151GAT : Nor_gate port map( I1 => G_6135GAT_OUT, I2 => G_6147GAT_OUT, O 
                           => G_6151GAT_OUT);
   G_6147GAT : Nor_gate port map( I1 => G_6124GAT_OUT, I2 => G_6141GAT_OUT, O 
                           => G_6147GAT_OUT);
   G_6146GAT : Inv_gate port map( I1 => G_6141GAT_OUT, O => G_6146GAT_OUT);
   G_6145GAT : Nor_gate port map( I1 => G_6138GAT_OUT, I2 => G_6141GAT_OUT, O 
                           => G_6145GAT_OUT);
   G_6141GAT : Inv_gate port map( I1 => G_6138GAT_OUT, O => G_6141GAT_OUT);
   G_6138GAT : Nor_gate port map( I1 => G_6133GAT_OUT, I2 => G_6134GAT_OUT, O 
                           => G_6138GAT_OUT);
   G_6135GAT : Nor_gate port map( I1 => G_6128GAT_OUT, I2 => G_6129GAT_OUT, O 
                           => G_6135GAT_OUT);
   G_6134GAT : Nor_gate port map( I1 => G_6124GAT_OUT, I2 => G_6108GAT_OUT, O 
                           => G_6134GAT_OUT);
   G_6133GAT : Nor_gate port map( I1 => G_6111GAT_OUT, I2 => G_6124GAT_OUT, O 
                           => G_6133GAT_OUT);
   G_6130GAT : Nor_gate port map( I1 => G_6118GAT_OUT, I2 => G_6119GAT_OUT, O 
                           => G_6130GAT_OUT);
   G_6129GAT : Nor_gate port map( I1 => G_6114GAT_OUT, I2 => G_6091GAT_OUT, O 
                           => G_6129GAT_OUT);
   G_6128GAT : Nor_gate port map( I1 => G_6094GAT_OUT, I2 => G_6114GAT_OUT, O 
                           => G_6128GAT_OUT);
   G_6124GAT : Nor_gate port map( I1 => G_6111GAT_OUT, I2 => G_6108GAT_OUT, O 
                           => G_6124GAT_OUT);
   G_6120GAT : Nor_gate port map( I1 => G_6101GAT_OUT, I2 => G_6102GAT_OUT, O 
                           => G_6120GAT_OUT);
   G_6119GAT : Nor_gate port map( I1 => G_6097GAT_OUT, I2 => G_6070GAT_OUT, O 
                           => G_6119GAT_OUT);
   G_6118GAT : Nor_gate port map( I1 => G_6073GAT_OUT, I2 => G_6097GAT_OUT, O 
                           => G_6118GAT_OUT);
   G_6114GAT : Nor_gate port map( I1 => G_6094GAT_OUT, I2 => G_6091GAT_OUT, O 
                           => G_6114GAT_OUT);
   G_6111GAT : Nor_gate port map( I1 => G_6089GAT_OUT, I2 => G_6090GAT_OUT, O 
                           => G_6111GAT_OUT);
   G_6108GAT : Nor_gate port map( I1 => G_6005GAT_OUT, I2 => G_6085GAT_OUT, O 
                           => G_6108GAT_OUT);
   G_6107GAT : Nor_gate port map( I1 => G_6085GAT_OUT, I2 => G_588GAT_OUT, O =>
                           G_6107GAT_OUT);
   G_6106GAT : Nor_gate port map( I1 => G_6061GAT_OUT, I2 => G_6085GAT_OUT, O 
                           => G_6106GAT_OUT);
   G_6103GAT : Nor_gate port map( I1 => G_6080GAT_OUT, I2 => G_6081GAT_OUT, O 
                           => G_6103GAT_OUT);
   G_6102GAT : Nor_gate port map( I1 => G_6076GAT_OUT, I2 => G_6046GAT_OUT, O 
                           => G_6102GAT_OUT);
   G_6101GAT : Nor_gate port map( I1 => G_6049GAT_OUT, I2 => G_6076GAT_OUT, O 
                           => G_6101GAT_OUT);
   G_6097GAT : Nor_gate port map( I1 => G_6073GAT_OUT, I2 => G_6070GAT_OUT, O 
                           => G_6097GAT_OUT);
   G_6094GAT : Nor_gate port map( I1 => G_6068GAT_OUT, I2 => G_6069GAT_OUT, O 
                           => G_6094GAT_OUT);
   G_6091GAT : Nor_gate port map( I1 => G_5975GAT_OUT, I2 => G_6064GAT_OUT, O 
                           => G_6091GAT_OUT);
   G_6090GAT : Nor_gate port map( I1 => G_6064GAT_OUT, I2 => G_636GAT_OUT, O =>
                           G_6090GAT_OUT);
   G_6089GAT : Nor_gate port map( I1 => G_6037GAT_OUT, I2 => G_6064GAT_OUT, O 
                           => G_6089GAT_OUT);
   G_6085GAT : Nor_gate port map( I1 => G_6061GAT_OUT, I2 => G_588GAT_OUT, O =>
                           G_6085GAT_OUT);
   G_6082GAT : Nor_gate port map( I1 => G_6056GAT_OUT, I2 => G_6057GAT_OUT, O 
                           => G_6082GAT_OUT);
   G_6081GAT : Nor_gate port map( I1 => G_6052GAT_OUT, I2 => G_6020GAT_OUT, O 
                           => G_6081GAT_OUT);
   G_6080GAT : Nor_gate port map( I1 => G_6023GAT_OUT, I2 => G_6052GAT_OUT, O 
                           => G_6080GAT_OUT);
   G_6076GAT : Nor_gate port map( I1 => G_6049GAT_OUT, I2 => G_6046GAT_OUT, O 
                           => G_6076GAT_OUT);
   G_6073GAT : Nor_gate port map( I1 => G_6044GAT_OUT, I2 => G_6045GAT_OUT, O 
                           => G_6073GAT_OUT);
   G_6070GAT : Nor_gate port map( I1 => G_5941GAT_OUT, I2 => G_6040GAT_OUT, O 
                           => G_6070GAT_OUT);
   G_6069GAT : Nor_gate port map( I1 => G_6040GAT_OUT, I2 => G_684GAT_OUT, O =>
                           G_6069GAT_OUT);
   G_6068GAT : Nor_gate port map( I1 => G_6011GAT_OUT, I2 => G_6040GAT_OUT, O 
                           => G_6068GAT_OUT);
   G_6064GAT : Nor_gate port map( I1 => G_6037GAT_OUT, I2 => G_636GAT_OUT, O =>
                           G_6064GAT_OUT);
   G_6061GAT : Nor_gate port map( I1 => G_6035GAT_OUT, I2 => G_6036GAT_OUT, O 
                           => G_6061GAT_OUT);
   G_6058GAT : Nor_gate port map( I1 => G_6030GAT_OUT, I2 => G_6031GAT_OUT, O 
                           => G_6058GAT_OUT);
   G_6057GAT : Nor_gate port map( I1 => G_6026GAT_OUT, I2 => G_5990GAT_OUT, O 
                           => G_6057GAT_OUT);
   G_6056GAT : Nor_gate port map( I1 => G_5993GAT_OUT, I2 => G_6026GAT_OUT, O 
                           => G_6056GAT_OUT);
   G_6052GAT : Nor_gate port map( I1 => G_6023GAT_OUT, I2 => G_6020GAT_OUT, O 
                           => G_6052GAT_OUT);
   G_6049GAT : Nor_gate port map( I1 => G_6018GAT_OUT, I2 => G_6019GAT_OUT, O 
                           => G_6049GAT_OUT);
   G_6046GAT : Nor_gate port map( I1 => G_5898GAT_OUT, I2 => G_6014GAT_OUT, O 
                           => G_6046GAT_OUT);
   G_6045GAT : Nor_gate port map( I1 => G_6014GAT_OUT, I2 => G_732GAT_OUT, O =>
                           G_6045GAT_OUT);
   G_6044GAT : Nor_gate port map( I1 => G_5981GAT_OUT, I2 => G_6014GAT_OUT, O 
                           => G_6044GAT_OUT);
   G_6040GAT : Nor_gate port map( I1 => G_6011GAT_OUT, I2 => G_684GAT_OUT, O =>
                           G_6040GAT_OUT);
   G_6037GAT : Nor_gate port map( I1 => G_6009GAT_OUT, I2 => G_6010GAT_OUT, O 
                           => G_6037GAT_OUT);
   G_6036GAT : Nor_gate port map( I1 => G_6005GAT_OUT, I2 => G_5930GAT_OUT, O 
                           => G_6036GAT_OUT);
   G_6035GAT : Nor_gate port map( I1 => G_5972GAT_OUT, I2 => G_6005GAT_OUT, O 
                           => G_6035GAT_OUT);
   G_6032GAT : Nor_gate port map( I1 => G_6000GAT_OUT, I2 => G_6001GAT_OUT, O 
                           => G_6032GAT_OUT);
   G_6031GAT : Nor_gate port map( I1 => G_5996GAT_OUT, I2 => G_5956GAT_OUT, O 
                           => G_6031GAT_OUT);
   G_6030GAT : Nor_gate port map( I1 => G_5959GAT_OUT, I2 => G_5996GAT_OUT, O 
                           => G_6030GAT_OUT);
   G_6026GAT : Nor_gate port map( I1 => G_5993GAT_OUT, I2 => G_5990GAT_OUT, O 
                           => G_6026GAT_OUT);
   G_6023GAT : Nor_gate port map( I1 => G_5988GAT_OUT, I2 => G_5989GAT_OUT, O 
                           => G_6023GAT_OUT);
   G_6020GAT : Nor_gate port map( I1 => G_5852GAT_OUT, I2 => G_5984GAT_OUT, O 
                           => G_6020GAT_OUT);
   G_6019GAT : Nor_gate port map( I1 => G_5984GAT_OUT, I2 => G_780GAT_OUT, O =>
                           G_6019GAT_OUT);
   G_6018GAT : Nor_gate port map( I1 => G_5947GAT_OUT, I2 => G_5984GAT_OUT, O 
                           => G_6018GAT_OUT);
   G_6014GAT : Nor_gate port map( I1 => G_5981GAT_OUT, I2 => G_732GAT_OUT, O =>
                           G_6014GAT_OUT);
   G_6011GAT : Nor_gate port map( I1 => G_5979GAT_OUT, I2 => G_5980GAT_OUT, O 
                           => G_6011GAT_OUT);
   G_6010GAT : Nor_gate port map( I1 => G_5975GAT_OUT, I2 => G_5935GAT_OUT, O 
                           => G_6010GAT_OUT);
   G_6009GAT : Nor_gate port map( I1 => G_5938GAT_OUT, I2 => G_5975GAT_OUT, O 
                           => G_6009GAT_OUT);
   G_6005GAT : Nor_gate port map( I1 => G_5972GAT_OUT, I2 => G_5930GAT_OUT, O 
                           => G_6005GAT_OUT);
   G_6002GAT : Nor_gate port map( I1 => G_5966GAT_OUT, I2 => G_5967GAT_OUT, O 
                           => G_6002GAT_OUT);
   G_6001GAT : Nor_gate port map( I1 => G_5962GAT_OUT, I2 => G_5913GAT_OUT, O 
                           => G_6001GAT_OUT);
   G_6000GAT : Nor_gate port map( I1 => G_5916GAT_OUT, I2 => G_5962GAT_OUT, O 
                           => G_6000GAT_OUT);
   G_5996GAT : Nor_gate port map( I1 => G_5959GAT_OUT, I2 => G_5956GAT_OUT, O 
                           => G_5996GAT_OUT);
   G_5993GAT : Nor_gate port map( I1 => G_5954GAT_OUT, I2 => G_5955GAT_OUT, O 
                           => G_5993GAT_OUT);
   G_5990GAT : Nor_gate port map( I1 => G_5804GAT_OUT, I2 => G_5950GAT_OUT, O 
                           => G_5990GAT_OUT);
   G_5989GAT : Nor_gate port map( I1 => G_5950GAT_OUT, I2 => G_828GAT_OUT, O =>
                           G_5989GAT_OUT);
   G_5988GAT : Nor_gate port map( I1 => G_5904GAT_OUT, I2 => G_5950GAT_OUT, O 
                           => G_5988GAT_OUT);
   G_5984GAT : Nor_gate port map( I1 => G_5947GAT_OUT, I2 => G_780GAT_OUT, O =>
                           G_5984GAT_OUT);
   G_5981GAT : Nor_gate port map( I1 => G_5945GAT_OUT, I2 => G_5946GAT_OUT, O 
                           => G_5981GAT_OUT);
   G_5980GAT : Nor_gate port map( I1 => G_5941GAT_OUT, I2 => G_5892GAT_OUT, O 
                           => G_5980GAT_OUT);
   G_5979GAT : Nor_gate port map( I1 => G_5895GAT_OUT, I2 => G_5941GAT_OUT, O 
                           => G_5979GAT_OUT);
   G_5975GAT : Nor_gate port map( I1 => G_5938GAT_OUT, I2 => G_5935GAT_OUT, O 
                           => G_5975GAT_OUT);
   G_5972GAT : Nor_gate port map( I1 => G_5933GAT_OUT, I2 => G_5934GAT_OUT, O 
                           => G_5972GAT_OUT);
   G_5968GAT : Nor_gate port map( I1 => G_5923GAT_OUT, I2 => G_5924GAT_OUT, O 
                           => G_5968GAT_OUT);
   G_5967GAT : Nor_gate port map( I1 => G_5919GAT_OUT, I2 => G_5867GAT_OUT, O 
                           => G_5967GAT_OUT);
   G_5966GAT : Nor_gate port map( I1 => G_5870GAT_OUT, I2 => G_5919GAT_OUT, O 
                           => G_5966GAT_OUT);
   G_5962GAT : Nor_gate port map( I1 => G_5916GAT_OUT, I2 => G_5913GAT_OUT, O 
                           => G_5962GAT_OUT);
   G_5959GAT : Nor_gate port map( I1 => G_5911GAT_OUT, I2 => G_5912GAT_OUT, O 
                           => G_5959GAT_OUT);
   G_5956GAT : Nor_gate port map( I1 => G_5755GAT_OUT, I2 => G_5907GAT_OUT, O 
                           => G_5956GAT_OUT);
   G_5955GAT : Nor_gate port map( I1 => G_5907GAT_OUT, I2 => G_876GAT_OUT, O =>
                           G_5955GAT_OUT);
   G_5954GAT : Nor_gate port map( I1 => G_5858GAT_OUT, I2 => G_5907GAT_OUT, O 
                           => G_5954GAT_OUT);
   G_5950GAT : Nor_gate port map( I1 => G_5904GAT_OUT, I2 => G_828GAT_OUT, O =>
                           G_5950GAT_OUT);
   G_5947GAT : Nor_gate port map( I1 => G_5902GAT_OUT, I2 => G_5903GAT_OUT, O 
                           => G_5947GAT_OUT);
   G_5946GAT : Nor_gate port map( I1 => G_5898GAT_OUT, I2 => G_5846GAT_OUT, O 
                           => G_5946GAT_OUT);
   G_5945GAT : Nor_gate port map( I1 => G_5849GAT_OUT, I2 => G_5898GAT_OUT, O 
                           => G_5945GAT_OUT);
   G_5941GAT : Nor_gate port map( I1 => G_5895GAT_OUT, I2 => G_5892GAT_OUT, O 
                           => G_5941GAT_OUT);
   G_5938GAT : Nor_gate port map( I1 => G_5890GAT_OUT, I2 => G_5891GAT_OUT, O 
                           => G_5938GAT_OUT);
   G_5935GAT : Nor_gate port map( I1 => G_5734GAT_OUT, I2 => G_5886GAT_OUT, O 
                           => G_5935GAT_OUT);
   G_5934GAT : Nor_gate port map( I1 => G_5886GAT_OUT, I2 => G_633GAT_OUT, O =>
                           G_5934GAT_OUT);
   G_5933GAT : Nor_gate port map( I1 => G_5837GAT_OUT, I2 => G_5886GAT_OUT, O 
                           => G_5933GAT_OUT);
   G_5930GAT : Nor_gate port map( I1 => G_5730GAT_OUT, I2 => G_5882GAT_OUT, O 
                           => G_5930GAT_OUT);
   G_5929GAT : Nor_gate port map( I1 => G_5882GAT_OUT, I2 => G_585GAT_OUT, O =>
                           G_5929GAT_OUT);
   G_5928GAT : Nor_gate port map( I1 => G_5834GAT_OUT, I2 => G_5882GAT_OUT, O 
                           => G_5928GAT_OUT);
   G_5925GAT : Nor_gate port map( I1 => G_5877GAT_OUT, I2 => G_5878GAT_OUT, O 
                           => G_5925GAT_OUT);
   G_5924GAT : Nor_gate port map( I1 => G_5873GAT_OUT, I2 => G_5819GAT_OUT, O 
                           => G_5924GAT_OUT);
   G_5923GAT : Nor_gate port map( I1 => G_5822GAT_OUT, I2 => G_5873GAT_OUT, O 
                           => G_5923GAT_OUT);
   G_5919GAT : Nor_gate port map( I1 => G_5870GAT_OUT, I2 => G_5867GAT_OUT, O 
                           => G_5919GAT_OUT);
   G_5916GAT : Nor_gate port map( I1 => G_5865GAT_OUT, I2 => G_5866GAT_OUT, O 
                           => G_5916GAT_OUT);
   G_5913GAT : Nor_gate port map( I1 => G_5700GAT_OUT, I2 => G_5861GAT_OUT, O 
                           => G_5913GAT_OUT);
   G_5912GAT : Nor_gate port map( I1 => G_5861GAT_OUT, I2 => G_924GAT_OUT, O =>
                           G_5912GAT_OUT);
   G_5911GAT : Nor_gate port map( I1 => G_5810GAT_OUT, I2 => G_5861GAT_OUT, O 
                           => G_5911GAT_OUT);
   G_5907GAT : Nor_gate port map( I1 => G_5858GAT_OUT, I2 => G_876GAT_OUT, O =>
                           G_5907GAT_OUT);
   G_5904GAT : Nor_gate port map( I1 => G_5856GAT_OUT, I2 => G_5857GAT_OUT, O 
                           => G_5904GAT_OUT);
   G_5903GAT : Nor_gate port map( I1 => G_5852GAT_OUT, I2 => G_5798GAT_OUT, O 
                           => G_5903GAT_OUT);
   G_5902GAT : Nor_gate port map( I1 => G_5801GAT_OUT, I2 => G_5852GAT_OUT, O 
                           => G_5902GAT_OUT);
   G_5898GAT : Nor_gate port map( I1 => G_5849GAT_OUT, I2 => G_5846GAT_OUT, O 
                           => G_5898GAT_OUT);
   G_5895GAT : Nor_gate port map( I1 => G_5844GAT_OUT, I2 => G_5845GAT_OUT, O 
                           => G_5895GAT_OUT);
   G_5892GAT : Nor_gate port map( I1 => G_5679GAT_OUT, I2 => G_5840GAT_OUT, O 
                           => G_5892GAT_OUT);
   G_5891GAT : Nor_gate port map( I1 => G_5840GAT_OUT, I2 => G_681GAT_OUT, O =>
                           G_5891GAT_OUT);
   G_5890GAT : Nor_gate port map( I1 => G_5789GAT_OUT, I2 => G_5840GAT_OUT, O 
                           => G_5890GAT_OUT);
   G_5886GAT : Nor_gate port map( I1 => G_5837GAT_OUT, I2 => G_633GAT_OUT, O =>
                           G_5886GAT_OUT);
   G_5882GAT : Nor_gate port map( I1 => G_5834GAT_OUT, I2 => G_585GAT_OUT, O =>
                           G_5882GAT_OUT);
   G_5879GAT : Nor_gate port map( I1 => G_5829GAT_OUT, I2 => G_5830GAT_OUT, O 
                           => G_5879GAT_OUT);
   G_5878GAT : Nor_gate port map( I1 => G_5825GAT_OUT, I2 => G_5770GAT_OUT, O 
                           => G_5878GAT_OUT);
   G_5877GAT : Nor_gate port map( I1 => G_5773GAT_OUT, I2 => G_5825GAT_OUT, O 
                           => G_5877GAT_OUT);
   G_5873GAT : Nor_gate port map( I1 => G_5822GAT_OUT, I2 => G_5819GAT_OUT, O 
                           => G_5873GAT_OUT);
   G_5870GAT : Nor_gate port map( I1 => G_5817GAT_OUT, I2 => G_5818GAT_OUT, O 
                           => G_5870GAT_OUT);
   G_5867GAT : Nor_gate port map( I1 => G_5645GAT_OUT, I2 => G_5813GAT_OUT, O 
                           => G_5867GAT_OUT);
   G_5866GAT : Nor_gate port map( I1 => G_5813GAT_OUT, I2 => G_972GAT_OUT, O =>
                           G_5866GAT_OUT);
   G_5865GAT : Nor_gate port map( I1 => G_5761GAT_OUT, I2 => G_5813GAT_OUT, O 
                           => G_5865GAT_OUT);
   G_5861GAT : Nor_gate port map( I1 => G_5810GAT_OUT, I2 => G_924GAT_OUT, O =>
                           G_5861GAT_OUT);
   G_5858GAT : Nor_gate port map( I1 => G_5808GAT_OUT, I2 => G_5809GAT_OUT, O 
                           => G_5858GAT_OUT);
   G_5857GAT : Nor_gate port map( I1 => G_5804GAT_OUT, I2 => G_5749GAT_OUT, O 
                           => G_5857GAT_OUT);
   G_5856GAT : Nor_gate port map( I1 => G_5752GAT_OUT, I2 => G_5804GAT_OUT, O 
                           => G_5856GAT_OUT);
   G_5852GAT : Nor_gate port map( I1 => G_5801GAT_OUT, I2 => G_5798GAT_OUT, O 
                           => G_5852GAT_OUT);
   G_5849GAT : Nor_gate port map( I1 => G_5796GAT_OUT, I2 => G_5797GAT_OUT, O 
                           => G_5849GAT_OUT);
   G_5846GAT : Nor_gate port map( I1 => G_5624GAT_OUT, I2 => G_5792GAT_OUT, O 
                           => G_5846GAT_OUT);
   G_5845GAT : Nor_gate port map( I1 => G_5792GAT_OUT, I2 => G_729GAT_OUT, O =>
                           G_5845GAT_OUT);
   G_5844GAT : Nor_gate port map( I1 => G_5740GAT_OUT, I2 => G_5792GAT_OUT, O 
                           => G_5844GAT_OUT);
   G_5840GAT : Nor_gate port map( I1 => G_5789GAT_OUT, I2 => G_681GAT_OUT, O =>
                           G_5840GAT_OUT);
   G_5837GAT : Nor_gate port map( I1 => G_5787GAT_OUT, I2 => G_5788GAT_OUT, O 
                           => G_5837GAT_OUT);
   G_5834GAT : Nor_gate port map( I1 => G_5785GAT_OUT, I2 => G_5786GAT_OUT, O 
                           => G_5834GAT_OUT);
   G_5831GAT : Nor_gate port map( I1 => G_5780GAT_OUT, I2 => G_5781GAT_OUT, O 
                           => G_5831GAT_OUT);
   G_5830GAT : Nor_gate port map( I1 => G_5776GAT_OUT, I2 => G_5715GAT_OUT, O 
                           => G_5830GAT_OUT);
   G_5829GAT : Nor_gate port map( I1 => G_5718GAT_OUT, I2 => G_5776GAT_OUT, O 
                           => G_5829GAT_OUT);
   G_5825GAT : Nor_gate port map( I1 => G_5773GAT_OUT, I2 => G_5770GAT_OUT, O 
                           => G_5825GAT_OUT);
   G_5822GAT : Nor_gate port map( I1 => G_5768GAT_OUT, I2 => G_5769GAT_OUT, O 
                           => G_5822GAT_OUT);
   G_5819GAT : Nor_gate port map( I1 => G_5581GAT_OUT, I2 => G_5764GAT_OUT, O 
                           => G_5819GAT_OUT);
   G_5818GAT : Nor_gate port map( I1 => G_5764GAT_OUT, I2 => G_1020GAT_OUT, O 
                           => G_5818GAT_OUT);
   G_5817GAT : Nor_gate port map( I1 => G_5706GAT_OUT, I2 => G_5764GAT_OUT, O 
                           => G_5817GAT_OUT);
   G_5813GAT : Nor_gate port map( I1 => G_5761GAT_OUT, I2 => G_972GAT_OUT, O =>
                           G_5813GAT_OUT);
   G_5810GAT : Nor_gate port map( I1 => G_5759GAT_OUT, I2 => G_5760GAT_OUT, O 
                           => G_5810GAT_OUT);
   G_5809GAT : Nor_gate port map( I1 => G_5755GAT_OUT, I2 => G_5694GAT_OUT, O 
                           => G_5809GAT_OUT);
   G_5808GAT : Nor_gate port map( I1 => G_5697GAT_OUT, I2 => G_5755GAT_OUT, O 
                           => G_5808GAT_OUT);
   G_5804GAT : Nor_gate port map( I1 => G_5752GAT_OUT, I2 => G_5749GAT_OUT, O 
                           => G_5804GAT_OUT);
   G_5801GAT : Nor_gate port map( I1 => G_5747GAT_OUT, I2 => G_5748GAT_OUT, O 
                           => G_5801GAT_OUT);
   G_5798GAT : Nor_gate port map( I1 => G_5560GAT_OUT, I2 => G_5743GAT_OUT, O 
                           => G_5798GAT_OUT);
   G_5797GAT : Nor_gate port map( I1 => G_5743GAT_OUT, I2 => G_777GAT_OUT, O =>
                           G_5797GAT_OUT);
   G_5796GAT : Nor_gate port map( I1 => G_5685GAT_OUT, I2 => G_5743GAT_OUT, O 
                           => G_5796GAT_OUT);
   G_5792GAT : Nor_gate port map( I1 => G_5740GAT_OUT, I2 => G_729GAT_OUT, O =>
                           G_5792GAT_OUT);
   G_5789GAT : Nor_gate port map( I1 => G_5738GAT_OUT, I2 => G_5739GAT_OUT, O 
                           => G_5789GAT_OUT);
   G_5788GAT : Nor_gate port map( I1 => G_5734GAT_OUT, I2 => G_5613GAT_OUT, O 
                           => G_5788GAT_OUT);
   G_5787GAT : Nor_gate port map( I1 => G_5676GAT_OUT, I2 => G_5734GAT_OUT, O 
                           => G_5787GAT_OUT);
   G_5786GAT : Nor_gate port map( I1 => G_5730GAT_OUT, I2 => G_5608GAT_OUT, O 
                           => G_5786GAT_OUT);
   G_5785GAT : Nor_gate port map( I1 => G_5673GAT_OUT, I2 => G_5730GAT_OUT, O 
                           => G_5785GAT_OUT);
   G_5782GAT : Nor_gate port map( I1 => G_5725GAT_OUT, I2 => G_5726GAT_OUT, O 
                           => G_5782GAT_OUT);
   G_5781GAT : Nor_gate port map( I1 => G_5721GAT_OUT, I2 => G_5660GAT_OUT, O 
                           => G_5781GAT_OUT);
   G_5780GAT : Nor_gate port map( I1 => G_5663GAT_OUT, I2 => G_5721GAT_OUT, O 
                           => G_5780GAT_OUT);
   G_5776GAT : Nor_gate port map( I1 => G_5718GAT_OUT, I2 => G_5715GAT_OUT, O 
                           => G_5776GAT_OUT);
   G_5773GAT : Nor_gate port map( I1 => G_5713GAT_OUT, I2 => G_5714GAT_OUT, O 
                           => G_5773GAT_OUT);
   G_5770GAT : Nor_gate port map( I1 => G_5522GAT_OUT, I2 => G_5709GAT_OUT, O 
                           => G_5770GAT_OUT);
   G_5769GAT : Nor_gate port map( I1 => G_5709GAT_OUT, I2 => G_1068GAT_OUT, O 
                           => G_5769GAT_OUT);
   G_5768GAT : Nor_gate port map( I1 => G_5651GAT_OUT, I2 => G_5709GAT_OUT, O 
                           => G_5768GAT_OUT);
   G_5764GAT : Nor_gate port map( I1 => G_5706GAT_OUT, I2 => G_1020GAT_OUT, O 
                           => G_5764GAT_OUT);
   G_5761GAT : Nor_gate port map( I1 => G_5704GAT_OUT, I2 => G_5705GAT_OUT, O 
                           => G_5761GAT_OUT);
   G_5760GAT : Nor_gate port map( I1 => G_5700GAT_OUT, I2 => G_5639GAT_OUT, O 
                           => G_5760GAT_OUT);
   G_5759GAT : Nor_gate port map( I1 => G_5642GAT_OUT, I2 => G_5700GAT_OUT, O 
                           => G_5759GAT_OUT);
   G_5755GAT : Nor_gate port map( I1 => G_5697GAT_OUT, I2 => G_5694GAT_OUT, O 
                           => G_5755GAT_OUT);
   G_5752GAT : Nor_gate port map( I1 => G_5692GAT_OUT, I2 => G_5693GAT_OUT, O 
                           => G_5752GAT_OUT);
   G_5749GAT : Nor_gate port map( I1 => G_5501GAT_OUT, I2 => G_5688GAT_OUT, O 
                           => G_5749GAT_OUT);
   G_5748GAT : Nor_gate port map( I1 => G_5688GAT_OUT, I2 => G_825GAT_OUT, O =>
                           G_5748GAT_OUT);
   G_5747GAT : Nor_gate port map( I1 => G_5630GAT_OUT, I2 => G_5688GAT_OUT, O 
                           => G_5747GAT_OUT);
   G_5743GAT : Nor_gate port map( I1 => G_5685GAT_OUT, I2 => G_777GAT_OUT, O =>
                           G_5743GAT_OUT);
   G_5740GAT : Nor_gate port map( I1 => G_5683GAT_OUT, I2 => G_5684GAT_OUT, O 
                           => G_5740GAT_OUT);
   G_5739GAT : Nor_gate port map( I1 => G_5679GAT_OUT, I2 => G_5618GAT_OUT, O 
                           => G_5739GAT_OUT);
   G_5738GAT : Nor_gate port map( I1 => G_5621GAT_OUT, I2 => G_5679GAT_OUT, O 
                           => G_5738GAT_OUT);
   G_5734GAT : Nor_gate port map( I1 => G_5676GAT_OUT, I2 => G_5613GAT_OUT, O 
                           => G_5734GAT_OUT);
   G_5730GAT : Nor_gate port map( I1 => G_5673GAT_OUT, I2 => G_5608GAT_OUT, O 
                           => G_5730GAT_OUT);
   G_5727GAT : Nor_gate port map( I1 => G_5670GAT_OUT, I2 => G_5671GAT_OUT, O 
                           => G_5727GAT_OUT);
   G_5726GAT : Nor_gate port map( I1 => G_5666GAT_OUT, I2 => G_5596GAT_OUT, O 
                           => G_5726GAT_OUT);
   G_5725GAT : Nor_gate port map( I1 => G_5599GAT_OUT, I2 => G_5666GAT_OUT, O 
                           => G_5725GAT_OUT);
   G_5721GAT : Nor_gate port map( I1 => G_5663GAT_OUT, I2 => G_5660GAT_OUT, O 
                           => G_5721GAT_OUT);
   G_5718GAT : Nor_gate port map( I1 => G_5658GAT_OUT, I2 => G_5659GAT_OUT, O 
                           => G_5718GAT_OUT);
   G_5715GAT : Nor_gate port map( I1 => G_5467GAT_OUT, I2 => G_5654GAT_OUT, O 
                           => G_5715GAT_OUT);
   G_5714GAT : Nor_gate port map( I1 => G_5654GAT_OUT, I2 => G_1116GAT_OUT, O 
                           => G_5714GAT_OUT);
   G_5713GAT : Nor_gate port map( I1 => G_5587GAT_OUT, I2 => G_5654GAT_OUT, O 
                           => G_5713GAT_OUT);
   G_5709GAT : Nor_gate port map( I1 => G_5651GAT_OUT, I2 => G_1068GAT_OUT, O 
                           => G_5709GAT_OUT);
   G_5706GAT : Nor_gate port map( I1 => G_5649GAT_OUT, I2 => G_5650GAT_OUT, O 
                           => G_5706GAT_OUT);
   G_5705GAT : Nor_gate port map( I1 => G_5645GAT_OUT, I2 => G_5575GAT_OUT, O 
                           => G_5705GAT_OUT);
   G_5704GAT : Nor_gate port map( I1 => G_5578GAT_OUT, I2 => G_5645GAT_OUT, O 
                           => G_5704GAT_OUT);
   G_5700GAT : Nor_gate port map( I1 => G_5642GAT_OUT, I2 => G_5639GAT_OUT, O 
                           => G_5700GAT_OUT);
   G_5697GAT : Nor_gate port map( I1 => G_5637GAT_OUT, I2 => G_5638GAT_OUT, O 
                           => G_5697GAT_OUT);
   G_5694GAT : Nor_gate port map( I1 => G_5446GAT_OUT, I2 => G_5633GAT_OUT, O 
                           => G_5694GAT_OUT);
   G_5693GAT : Nor_gate port map( I1 => G_5633GAT_OUT, I2 => G_873GAT_OUT, O =>
                           G_5693GAT_OUT);
   G_5692GAT : Nor_gate port map( I1 => G_5566GAT_OUT, I2 => G_5633GAT_OUT, O 
                           => G_5692GAT_OUT);
   G_5688GAT : Nor_gate port map( I1 => G_5630GAT_OUT, I2 => G_825GAT_OUT, O =>
                           G_5688GAT_OUT);
   G_5685GAT : Nor_gate port map( I1 => G_5628GAT_OUT, I2 => G_5629GAT_OUT, O 
                           => G_5685GAT_OUT);
   G_5684GAT : Nor_gate port map( I1 => G_5624GAT_OUT, I2 => G_5554GAT_OUT, O 
                           => G_5684GAT_OUT);
   G_5683GAT : Nor_gate port map( I1 => G_5557GAT_OUT, I2 => G_5624GAT_OUT, O 
                           => G_5683GAT_OUT);
   G_5679GAT : Nor_gate port map( I1 => G_5621GAT_OUT, I2 => G_5618GAT_OUT, O 
                           => G_5679GAT_OUT);
   G_5676GAT : Nor_gate port map( I1 => G_5616GAT_OUT, I2 => G_5617GAT_OUT, O 
                           => G_5676GAT_OUT);
   G_5673GAT : Nor_gate port map( I1 => G_5611GAT_OUT, I2 => G_5612GAT_OUT, O 
                           => G_5673GAT_OUT);
   G_5671GAT : Nor_gate port map( I1 => G_5602GAT_OUT, I2 => G_5537GAT_OUT, O 
                           => G_5671GAT_OUT);
   G_5670GAT : Nor_gate port map( I1 => G_1308GAT_OUT, I2 => G_5602GAT_OUT, O 
                           => G_5670GAT_OUT);
   G_5666GAT : Nor_gate port map( I1 => G_5599GAT_OUT, I2 => G_5596GAT_OUT, O 
                           => G_5666GAT_OUT);
   G_5663GAT : Nor_gate port map( I1 => G_5594GAT_OUT, I2 => G_5595GAT_OUT, O 
                           => G_5663GAT_OUT);
   G_5660GAT : Nor_gate port map( I1 => G_5416GAT_OUT, I2 => G_5590GAT_OUT, O 
                           => G_5660GAT_OUT);
   G_5659GAT : Nor_gate port map( I1 => G_5590GAT_OUT, I2 => G_1164GAT_OUT, O 
                           => G_5659GAT_OUT);
   G_5658GAT : Nor_gate port map( I1 => G_5528GAT_OUT, I2 => G_5590GAT_OUT, O 
                           => G_5658GAT_OUT);
   G_5654GAT : Nor_gate port map( I1 => G_5587GAT_OUT, I2 => G_1116GAT_OUT, O 
                           => G_5654GAT_OUT);
   G_5651GAT : Nor_gate port map( I1 => G_5585GAT_OUT, I2 => G_5586GAT_OUT, O 
                           => G_5651GAT_OUT);
   G_5650GAT : Nor_gate port map( I1 => G_5581GAT_OUT, I2 => G_5516GAT_OUT, O 
                           => G_5650GAT_OUT);
   G_5649GAT : Nor_gate port map( I1 => G_5519GAT_OUT, I2 => G_5581GAT_OUT, O 
                           => G_5649GAT_OUT);
   G_5645GAT : Nor_gate port map( I1 => G_5578GAT_OUT, I2 => G_5575GAT_OUT, O 
                           => G_5645GAT_OUT);
   G_5642GAT : Nor_gate port map( I1 => G_5573GAT_OUT, I2 => G_5574GAT_OUT, O 
                           => G_5642GAT_OUT);
   G_5639GAT : Nor_gate port map( I1 => G_5395GAT_OUT, I2 => G_5569GAT_OUT, O 
                           => G_5639GAT_OUT);
   G_5638GAT : Nor_gate port map( I1 => G_5569GAT_OUT, I2 => G_921GAT_OUT, O =>
                           G_5638GAT_OUT);
   G_5637GAT : Nor_gate port map( I1 => G_5507GAT_OUT, I2 => G_5569GAT_OUT, O 
                           => G_5637GAT_OUT);
   G_5633GAT : Nor_gate port map( I1 => G_5566GAT_OUT, I2 => G_873GAT_OUT, O =>
                           G_5633GAT_OUT);
   G_5630GAT : Nor_gate port map( I1 => G_5564GAT_OUT, I2 => G_5565GAT_OUT, O 
                           => G_5630GAT_OUT);
   G_5629GAT : Nor_gate port map( I1 => G_5560GAT_OUT, I2 => G_5495GAT_OUT, O 
                           => G_5629GAT_OUT);
   G_5628GAT : Nor_gate port map( I1 => G_5498GAT_OUT, I2 => G_5560GAT_OUT, O 
                           => G_5628GAT_OUT);
   G_5624GAT : Nor_gate port map( I1 => G_5557GAT_OUT, I2 => G_5554GAT_OUT, O 
                           => G_5624GAT_OUT);
   G_5621GAT : Nor_gate port map( I1 => G_5552GAT_OUT, I2 => G_5553GAT_OUT, O 
                           => G_5621GAT_OUT);
   G_5618GAT : Nor_gate port map( I1 => G_5374GAT_OUT, I2 => G_5548GAT_OUT, O 
                           => G_5618GAT_OUT);
   G_5617GAT : Nor_gate port map( I1 => G_5548GAT_OUT, I2 => G_678GAT_OUT, O =>
                           G_5617GAT_OUT);
   G_5616GAT : Nor_gate port map( I1 => G_5486GAT_OUT, I2 => G_5548GAT_OUT, O 
                           => G_5616GAT_OUT);
   G_5613GAT : Nor_gate port map( I1 => G_5370GAT_OUT, I2 => G_5544GAT_OUT, O 
                           => G_5613GAT_OUT);
   G_5612GAT : Nor_gate port map( I1 => G_5544GAT_OUT, I2 => G_630GAT_OUT, O =>
                           G_5612GAT_OUT);
   G_5611GAT : Nor_gate port map( I1 => G_5483GAT_OUT, I2 => G_5544GAT_OUT, O 
                           => G_5611GAT_OUT);
   G_5608GAT : Nor_gate port map( I1 => G_5366GAT_OUT, I2 => G_5540GAT_OUT, O 
                           => G_5608GAT_OUT);
   G_5607GAT : Nor_gate port map( I1 => G_5540GAT_OUT, I2 => G_582GAT_OUT, O =>
                           G_5607GAT_OUT);
   G_5606GAT : Nor_gate port map( I1 => G_5480GAT_OUT, I2 => G_5540GAT_OUT, O 
                           => G_5606GAT_OUT);
   G_5602GAT : Nor_gate port map( I1 => G_1308GAT_OUT, I2 => G_5537GAT_OUT, O 
                           => G_5602GAT_OUT);
   G_5599GAT : Nor_gate port map( I1 => G_5535GAT_OUT, I2 => G_5536GAT_OUT, O 
                           => G_5599GAT_OUT);
   G_5596GAT : Nor_gate port map( I1 => G_5360GAT_OUT, I2 => G_5531GAT_OUT, O 
                           => G_5596GAT_OUT);
   G_5595GAT : Nor_gate port map( I1 => G_5531GAT_OUT, I2 => G_1212GAT_OUT, O 
                           => G_5595GAT_OUT);
   G_5594GAT : Nor_gate port map( I1 => G_5473GAT_OUT, I2 => G_5531GAT_OUT, O 
                           => G_5594GAT_OUT);
   G_5590GAT : Nor_gate port map( I1 => G_5528GAT_OUT, I2 => G_1164GAT_OUT, O 
                           => G_5590GAT_OUT);
   G_5587GAT : Nor_gate port map( I1 => G_5526GAT_OUT, I2 => G_5527GAT_OUT, O 
                           => G_5587GAT_OUT);
   G_5586GAT : Nor_gate port map( I1 => G_5522GAT_OUT, I2 => G_5461GAT_OUT, O 
                           => G_5586GAT_OUT);
   G_5585GAT : Nor_gate port map( I1 => G_5464GAT_OUT, I2 => G_5522GAT_OUT, O 
                           => G_5585GAT_OUT);
   G_5581GAT : Nor_gate port map( I1 => G_5519GAT_OUT, I2 => G_5516GAT_OUT, O 
                           => G_5581GAT_OUT);
   G_5578GAT : Nor_gate port map( I1 => G_5514GAT_OUT, I2 => G_5515GAT_OUT, O 
                           => G_5578GAT_OUT);
   G_5575GAT : Nor_gate port map( I1 => G_5339GAT_OUT, I2 => G_5510GAT_OUT, O 
                           => G_5575GAT_OUT);
   G_5574GAT : Nor_gate port map( I1 => G_5510GAT_OUT, I2 => G_969GAT_OUT, O =>
                           G_5574GAT_OUT);
   G_5573GAT : Nor_gate port map( I1 => G_5452GAT_OUT, I2 => G_5510GAT_OUT, O 
                           => G_5573GAT_OUT);
   G_5569GAT : Nor_gate port map( I1 => G_5507GAT_OUT, I2 => G_921GAT_OUT, O =>
                           G_5569GAT_OUT);
   G_5566GAT : Nor_gate port map( I1 => G_5505GAT_OUT, I2 => G_5506GAT_OUT, O 
                           => G_5566GAT_OUT);
   G_5565GAT : Nor_gate port map( I1 => G_5501GAT_OUT, I2 => G_5440GAT_OUT, O 
                           => G_5565GAT_OUT);
   G_5564GAT : Nor_gate port map( I1 => G_5443GAT_OUT, I2 => G_5501GAT_OUT, O 
                           => G_5564GAT_OUT);
   G_5560GAT : Nor_gate port map( I1 => G_5498GAT_OUT, I2 => G_5495GAT_OUT, O 
                           => G_5560GAT_OUT);
   G_5557GAT : Nor_gate port map( I1 => G_5493GAT_OUT, I2 => G_5494GAT_OUT, O 
                           => G_5557GAT_OUT);
   G_5554GAT : Nor_gate port map( I1 => G_5318GAT_OUT, I2 => G_5489GAT_OUT, O 
                           => G_5554GAT_OUT);
   G_5553GAT : Nor_gate port map( I1 => G_5489GAT_OUT, I2 => G_726GAT_OUT, O =>
                           G_5553GAT_OUT);
   G_5552GAT : Nor_gate port map( I1 => G_5431GAT_OUT, I2 => G_5489GAT_OUT, O 
                           => G_5552GAT_OUT);
   G_5548GAT : Nor_gate port map( I1 => G_5486GAT_OUT, I2 => G_678GAT_OUT, O =>
                           G_5548GAT_OUT);
   G_5544GAT : Nor_gate port map( I1 => G_5483GAT_OUT, I2 => G_630GAT_OUT, O =>
                           G_5544GAT_OUT);
   G_5540GAT : Nor_gate port map( I1 => G_5480GAT_OUT, I2 => G_582GAT_OUT, O =>
                           G_5540GAT_OUT);
   G_5537GAT : Nor_gate port map( I1 => G_5304GAT_OUT, I2 => G_5476GAT_OUT, O 
                           => G_5537GAT_OUT);
   G_5536GAT : Nor_gate port map( I1 => G_5476GAT_OUT, I2 => G_1260GAT_OUT, O 
                           => G_5536GAT_OUT);
   G_5535GAT : Nor_gate port map( I1 => G_5422GAT_OUT, I2 => G_5476GAT_OUT, O 
                           => G_5535GAT_OUT);
   G_5531GAT : Nor_gate port map( I1 => G_5473GAT_OUT, I2 => G_1212GAT_OUT, O 
                           => G_5531GAT_OUT);
   G_5528GAT : Nor_gate port map( I1 => G_5471GAT_OUT, I2 => G_5472GAT_OUT, O 
                           => G_5528GAT_OUT);
   G_5527GAT : Nor_gate port map( I1 => G_5467GAT_OUT, I2 => G_5410GAT_OUT, O 
                           => G_5527GAT_OUT);
   G_5526GAT : Nor_gate port map( I1 => G_5413GAT_OUT, I2 => G_5467GAT_OUT, O 
                           => G_5526GAT_OUT);
   G_5522GAT : Nor_gate port map( I1 => G_5464GAT_OUT, I2 => G_5461GAT_OUT, O 
                           => G_5522GAT_OUT);
   G_5519GAT : Nor_gate port map( I1 => G_5459GAT_OUT, I2 => G_5460GAT_OUT, O 
                           => G_5519GAT_OUT);
   G_5516GAT : Nor_gate port map( I1 => G_5283GAT_OUT, I2 => G_5455GAT_OUT, O 
                           => G_5516GAT_OUT);
   G_5515GAT : Nor_gate port map( I1 => G_5455GAT_OUT, I2 => G_1017GAT_OUT, O 
                           => G_5515GAT_OUT);
   G_5514GAT : Nor_gate port map( I1 => G_5401GAT_OUT, I2 => G_5455GAT_OUT, O 
                           => G_5514GAT_OUT);
   G_5510GAT : Nor_gate port map( I1 => G_5452GAT_OUT, I2 => G_969GAT_OUT, O =>
                           G_5510GAT_OUT);
   G_5507GAT : Nor_gate port map( I1 => G_5450GAT_OUT, I2 => G_5451GAT_OUT, O 
                           => G_5507GAT_OUT);
   G_5506GAT : Nor_gate port map( I1 => G_5446GAT_OUT, I2 => G_5389GAT_OUT, O 
                           => G_5506GAT_OUT);
   G_5505GAT : Nor_gate port map( I1 => G_5392GAT_OUT, I2 => G_5446GAT_OUT, O 
                           => G_5505GAT_OUT);
   G_5501GAT : Nor_gate port map( I1 => G_5443GAT_OUT, I2 => G_5440GAT_OUT, O 
                           => G_5501GAT_OUT);
   G_5498GAT : Nor_gate port map( I1 => G_5438GAT_OUT, I2 => G_5439GAT_OUT, O 
                           => G_5498GAT_OUT);
   G_5495GAT : Nor_gate port map( I1 => G_5262GAT_OUT, I2 => G_5434GAT_OUT, O 
                           => G_5495GAT_OUT);
   G_5494GAT : Nor_gate port map( I1 => G_5434GAT_OUT, I2 => G_774GAT_OUT, O =>
                           G_5494GAT_OUT);
   G_5493GAT : Nor_gate port map( I1 => G_5380GAT_OUT, I2 => G_5434GAT_OUT, O 
                           => G_5493GAT_OUT);
   G_5489GAT : Nor_gate port map( I1 => G_5431GAT_OUT, I2 => G_726GAT_OUT, O =>
                           G_5489GAT_OUT);
   G_5486GAT : Nor_gate port map( I1 => G_5429GAT_OUT, I2 => G_5430GAT_OUT, O 
                           => G_5486GAT_OUT);
   G_5483GAT : Nor_gate port map( I1 => G_5427GAT_OUT, I2 => G_5428GAT_OUT, O 
                           => G_5483GAT_OUT);
   G_5480GAT : Nor_gate port map( I1 => G_5425GAT_OUT, I2 => G_5426GAT_OUT, O 
                           => G_5480GAT_OUT);
   G_5476GAT : Nor_gate port map( I1 => G_5422GAT_OUT, I2 => G_1260GAT_OUT, O 
                           => G_5476GAT_OUT);
   G_5473GAT : Nor_gate port map( I1 => G_5420GAT_OUT, I2 => G_5421GAT_OUT, O 
                           => G_5473GAT_OUT);
   G_5472GAT : Nor_gate port map( I1 => G_5416GAT_OUT, I2 => G_5354GAT_OUT, O 
                           => G_5472GAT_OUT);
   G_5471GAT : Nor_gate port map( I1 => G_5357GAT_OUT, I2 => G_5416GAT_OUT, O 
                           => G_5471GAT_OUT);
   G_5467GAT : Nor_gate port map( I1 => G_5413GAT_OUT, I2 => G_5410GAT_OUT, O 
                           => G_5467GAT_OUT);
   G_5464GAT : Nor_gate port map( I1 => G_5408GAT_OUT, I2 => G_5409GAT_OUT, O 
                           => G_5464GAT_OUT);
   G_5461GAT : Nor_gate port map( I1 => G_5221GAT_OUT, I2 => G_5404GAT_OUT, O 
                           => G_5461GAT_OUT);
   G_5460GAT : Nor_gate port map( I1 => G_5404GAT_OUT, I2 => G_1065GAT_OUT, O 
                           => G_5460GAT_OUT);
   G_5459GAT : Nor_gate port map( I1 => G_5345GAT_OUT, I2 => G_5404GAT_OUT, O 
                           => G_5459GAT_OUT);
   G_5455GAT : Nor_gate port map( I1 => G_5401GAT_OUT, I2 => G_1017GAT_OUT, O 
                           => G_5455GAT_OUT);
   G_5452GAT : Nor_gate port map( I1 => G_5399GAT_OUT, I2 => G_5400GAT_OUT, O 
                           => G_5452GAT_OUT);
   G_5451GAT : Nor_gate port map( I1 => G_5395GAT_OUT, I2 => G_5333GAT_OUT, O 
                           => G_5451GAT_OUT);
   G_5450GAT : Nor_gate port map( I1 => G_5336GAT_OUT, I2 => G_5395GAT_OUT, O 
                           => G_5450GAT_OUT);
   G_5446GAT : Nor_gate port map( I1 => G_5392GAT_OUT, I2 => G_5389GAT_OUT, O 
                           => G_5446GAT_OUT);
   G_5443GAT : Nor_gate port map( I1 => G_5387GAT_OUT, I2 => G_5388GAT_OUT, O 
                           => G_5443GAT_OUT);
   G_5440GAT : Nor_gate port map( I1 => G_5200GAT_OUT, I2 => G_5383GAT_OUT, O 
                           => G_5440GAT_OUT);
   G_5439GAT : Nor_gate port map( I1 => G_5383GAT_OUT, I2 => G_822GAT_OUT, O =>
                           G_5439GAT_OUT);
   G_5438GAT : Nor_gate port map( I1 => G_5324GAT_OUT, I2 => G_5383GAT_OUT, O 
                           => G_5438GAT_OUT);
   G_5434GAT : Nor_gate port map( I1 => G_5380GAT_OUT, I2 => G_774GAT_OUT, O =>
                           G_5434GAT_OUT);
   G_5431GAT : Nor_gate port map( I1 => G_5378GAT_OUT, I2 => G_5379GAT_OUT, O 
                           => G_5431GAT_OUT);
   G_5430GAT : Nor_gate port map( I1 => G_5374GAT_OUT, I2 => G_5251GAT_OUT, O 
                           => G_5430GAT_OUT);
   G_5429GAT : Nor_gate port map( I1 => G_5315GAT_OUT, I2 => G_5374GAT_OUT, O 
                           => G_5429GAT_OUT);
   G_5428GAT : Nor_gate port map( I1 => G_5370GAT_OUT, I2 => G_5246GAT_OUT, O 
                           => G_5428GAT_OUT);
   G_5427GAT : Nor_gate port map( I1 => G_5312GAT_OUT, I2 => G_5370GAT_OUT, O 
                           => G_5427GAT_OUT);
   G_5426GAT : Nor_gate port map( I1 => G_5366GAT_OUT, I2 => G_5241GAT_OUT, O 
                           => G_5426GAT_OUT);
   G_5425GAT : Nor_gate port map( I1 => G_5309GAT_OUT, I2 => G_5366GAT_OUT, O 
                           => G_5425GAT_OUT);
   G_5422GAT : Nor_gate port map( I1 => G_5364GAT_OUT, I2 => G_5365GAT_OUT, O 
                           => G_5422GAT_OUT);
   G_5421GAT : Nor_gate port map( I1 => G_5360GAT_OUT, I2 => G_5298GAT_OUT, O 
                           => G_5421GAT_OUT);
   G_5420GAT : Nor_gate port map( I1 => G_5301GAT_OUT, I2 => G_5360GAT_OUT, O 
                           => G_5420GAT_OUT);
   G_5416GAT : Nor_gate port map( I1 => G_5357GAT_OUT, I2 => G_5354GAT_OUT, O 
                           => G_5416GAT_OUT);
   G_5413GAT : Nor_gate port map( I1 => G_5352GAT_OUT, I2 => G_5353GAT_OUT, O 
                           => G_5413GAT_OUT);
   G_5410GAT : Nor_gate port map( I1 => G_5163GAT_OUT, I2 => G_5348GAT_OUT, O 
                           => G_5410GAT_OUT);
   G_5409GAT : Nor_gate port map( I1 => G_5348GAT_OUT, I2 => G_1113GAT_OUT, O 
                           => G_5409GAT_OUT);
   G_5408GAT : Nor_gate port map( I1 => G_5289GAT_OUT, I2 => G_5348GAT_OUT, O 
                           => G_5408GAT_OUT);
   G_5404GAT : Nor_gate port map( I1 => G_5345GAT_OUT, I2 => G_1065GAT_OUT, O 
                           => G_5404GAT_OUT);
   G_5401GAT : Nor_gate port map( I1 => G_5343GAT_OUT, I2 => G_5344GAT_OUT, O 
                           => G_5401GAT_OUT);
   G_5400GAT : Nor_gate port map( I1 => G_5339GAT_OUT, I2 => G_5277GAT_OUT, O 
                           => G_5400GAT_OUT);
   G_5399GAT : Nor_gate port map( I1 => G_5280GAT_OUT, I2 => G_5339GAT_OUT, O 
                           => G_5399GAT_OUT);
   G_5395GAT : Nor_gate port map( I1 => G_5336GAT_OUT, I2 => G_5333GAT_OUT, O 
                           => G_5395GAT_OUT);
   G_5392GAT : Nor_gate port map( I1 => G_5331GAT_OUT, I2 => G_5332GAT_OUT, O 
                           => G_5392GAT_OUT);
   G_5389GAT : Nor_gate port map( I1 => G_5142GAT_OUT, I2 => G_5327GAT_OUT, O 
                           => G_5389GAT_OUT);
   G_5388GAT : Nor_gate port map( I1 => G_5327GAT_OUT, I2 => G_870GAT_OUT, O =>
                           G_5388GAT_OUT);
   G_5387GAT : Nor_gate port map( I1 => G_5268GAT_OUT, I2 => G_5327GAT_OUT, O 
                           => G_5387GAT_OUT);
   G_5383GAT : Nor_gate port map( I1 => G_5324GAT_OUT, I2 => G_822GAT_OUT, O =>
                           G_5383GAT_OUT);
   G_5380GAT : Nor_gate port map( I1 => G_5322GAT_OUT, I2 => G_5323GAT_OUT, O 
                           => G_5380GAT_OUT);
   G_5379GAT : Nor_gate port map( I1 => G_5318GAT_OUT, I2 => G_5256GAT_OUT, O 
                           => G_5379GAT_OUT);
   G_5378GAT : Nor_gate port map( I1 => G_5259GAT_OUT, I2 => G_5318GAT_OUT, O 
                           => G_5378GAT_OUT);
   G_5374GAT : Nor_gate port map( I1 => G_5315GAT_OUT, I2 => G_5251GAT_OUT, O 
                           => G_5374GAT_OUT);
   G_5370GAT : Nor_gate port map( I1 => G_5312GAT_OUT, I2 => G_5246GAT_OUT, O 
                           => G_5370GAT_OUT);
   G_5366GAT : Nor_gate port map( I1 => G_5309GAT_OUT, I2 => G_5241GAT_OUT, O 
                           => G_5366GAT_OUT);
   G_5365GAT : Nor_gate port map( I1 => G_5304GAT_OUT, I2 => G_5236GAT_OUT, O 
                           => G_5365GAT_OUT);
   G_5364GAT : Nor_gate port map( I1 => G_1305GAT_OUT, I2 => G_5304GAT_OUT, O 
                           => G_5364GAT_OUT);
   G_5360GAT : Nor_gate port map( I1 => G_5301GAT_OUT, I2 => G_5298GAT_OUT, O 
                           => G_5360GAT_OUT);
   G_5357GAT : Nor_gate port map( I1 => G_5296GAT_OUT, I2 => G_5297GAT_OUT, O 
                           => G_5357GAT_OUT);
   G_5354GAT : Nor_gate port map( I1 => G_5109GAT_OUT, I2 => G_5292GAT_OUT, O 
                           => G_5354GAT_OUT);
   G_5353GAT : Nor_gate port map( I1 => G_5292GAT_OUT, I2 => G_1161GAT_OUT, O 
                           => G_5353GAT_OUT);
   G_5352GAT : Nor_gate port map( I1 => G_5227GAT_OUT, I2 => G_5292GAT_OUT, O 
                           => G_5352GAT_OUT);
   G_5348GAT : Nor_gate port map( I1 => G_5289GAT_OUT, I2 => G_1113GAT_OUT, O 
                           => G_5348GAT_OUT);
   G_5345GAT : Nor_gate port map( I1 => G_5287GAT_OUT, I2 => G_5288GAT_OUT, O 
                           => G_5345GAT_OUT);
   G_5344GAT : Nor_gate port map( I1 => G_5283GAT_OUT, I2 => G_5215GAT_OUT, O 
                           => G_5344GAT_OUT);
   G_5343GAT : Nor_gate port map( I1 => G_5218GAT_OUT, I2 => G_5283GAT_OUT, O 
                           => G_5343GAT_OUT);
   G_5339GAT : Nor_gate port map( I1 => G_5280GAT_OUT, I2 => G_5277GAT_OUT, O 
                           => G_5339GAT_OUT);
   G_5336GAT : Nor_gate port map( I1 => G_5275GAT_OUT, I2 => G_5276GAT_OUT, O 
                           => G_5336GAT_OUT);
   G_5333GAT : Nor_gate port map( I1 => G_5088GAT_OUT, I2 => G_5271GAT_OUT, O 
                           => G_5333GAT_OUT);
   G_5332GAT : Nor_gate port map( I1 => G_5271GAT_OUT, I2 => G_918GAT_OUT, O =>
                           G_5332GAT_OUT);
   G_5331GAT : Nor_gate port map( I1 => G_5206GAT_OUT, I2 => G_5271GAT_OUT, O 
                           => G_5331GAT_OUT);
   G_5327GAT : Nor_gate port map( I1 => G_5268GAT_OUT, I2 => G_870GAT_OUT, O =>
                           G_5327GAT_OUT);
   G_5324GAT : Nor_gate port map( I1 => G_5266GAT_OUT, I2 => G_5267GAT_OUT, O 
                           => G_5324GAT_OUT);
   G_5323GAT : Nor_gate port map( I1 => G_5262GAT_OUT, I2 => G_5194GAT_OUT, O 
                           => G_5323GAT_OUT);
   G_5322GAT : Nor_gate port map( I1 => G_5197GAT_OUT, I2 => G_5262GAT_OUT, O 
                           => G_5322GAT_OUT);
   G_5318GAT : Nor_gate port map( I1 => G_5259GAT_OUT, I2 => G_5256GAT_OUT, O 
                           => G_5318GAT_OUT);
   G_5315GAT : Nor_gate port map( I1 => G_5254GAT_OUT, I2 => G_5255GAT_OUT, O 
                           => G_5315GAT_OUT);
   G_5312GAT : Nor_gate port map( I1 => G_5249GAT_OUT, I2 => G_5250GAT_OUT, O 
                           => G_5312GAT_OUT);
   G_5309GAT : Nor_gate port map( I1 => G_5244GAT_OUT, I2 => G_5245GAT_OUT, O 
                           => G_5309GAT_OUT);
   G_5304GAT : Nor_gate port map( I1 => G_1305GAT_OUT, I2 => G_5236GAT_OUT, O 
                           => G_5304GAT_OUT);
   G_5301GAT : Nor_gate port map( I1 => G_5234GAT_OUT, I2 => G_5235GAT_OUT, O 
                           => G_5301GAT_OUT);
   G_5298GAT : Nor_gate port map( I1 => G_5059GAT_OUT, I2 => G_5230GAT_OUT, O 
                           => G_5298GAT_OUT);
   G_5297GAT : Nor_gate port map( I1 => G_5230GAT_OUT, I2 => G_1209GAT_OUT, O 
                           => G_5297GAT_OUT);
   G_5296GAT : Nor_gate port map( I1 => G_5169GAT_OUT, I2 => G_5230GAT_OUT, O 
                           => G_5296GAT_OUT);
   G_5292GAT : Nor_gate port map( I1 => G_5227GAT_OUT, I2 => G_1161GAT_OUT, O 
                           => G_5292GAT_OUT);
   G_5289GAT : Nor_gate port map( I1 => G_5225GAT_OUT, I2 => G_5226GAT_OUT, O 
                           => G_5289GAT_OUT);
   G_5288GAT : Nor_gate port map( I1 => G_5221GAT_OUT, I2 => G_5157GAT_OUT, O 
                           => G_5288GAT_OUT);
   G_5287GAT : Nor_gate port map( I1 => G_5160GAT_OUT, I2 => G_5221GAT_OUT, O 
                           => G_5287GAT_OUT);
   G_5283GAT : Nor_gate port map( I1 => G_5218GAT_OUT, I2 => G_5215GAT_OUT, O 
                           => G_5283GAT_OUT);
   G_5280GAT : Nor_gate port map( I1 => G_5213GAT_OUT, I2 => G_5214GAT_OUT, O 
                           => G_5280GAT_OUT);
   G_5277GAT : Nor_gate port map( I1 => G_5038GAT_OUT, I2 => G_5209GAT_OUT, O 
                           => G_5277GAT_OUT);
   G_5276GAT : Nor_gate port map( I1 => G_5209GAT_OUT, I2 => G_966GAT_OUT, O =>
                           G_5276GAT_OUT);
   G_5275GAT : Nor_gate port map( I1 => G_5148GAT_OUT, I2 => G_5209GAT_OUT, O 
                           => G_5275GAT_OUT);
   G_5271GAT : Nor_gate port map( I1 => G_5206GAT_OUT, I2 => G_918GAT_OUT, O =>
                           G_5271GAT_OUT);
   G_5268GAT : Nor_gate port map( I1 => G_5204GAT_OUT, I2 => G_5205GAT_OUT, O 
                           => G_5268GAT_OUT);
   G_5267GAT : Nor_gate port map( I1 => G_5200GAT_OUT, I2 => G_5136GAT_OUT, O 
                           => G_5267GAT_OUT);
   G_5266GAT : Nor_gate port map( I1 => G_5139GAT_OUT, I2 => G_5200GAT_OUT, O 
                           => G_5266GAT_OUT);
   G_5262GAT : Nor_gate port map( I1 => G_5197GAT_OUT, I2 => G_5194GAT_OUT, O 
                           => G_5262GAT_OUT);
   G_5259GAT : Nor_gate port map( I1 => G_5192GAT_OUT, I2 => G_5193GAT_OUT, O 
                           => G_5259GAT_OUT);
   G_5256GAT : Nor_gate port map( I1 => G_5017GAT_OUT, I2 => G_5188GAT_OUT, O 
                           => G_5256GAT_OUT);
   G_5255GAT : Nor_gate port map( I1 => G_5188GAT_OUT, I2 => G_723GAT_OUT, O =>
                           G_5255GAT_OUT);
   G_5254GAT : Nor_gate port map( I1 => G_5127GAT_OUT, I2 => G_5188GAT_OUT, O 
                           => G_5254GAT_OUT);
   G_5251GAT : Nor_gate port map( I1 => G_5013GAT_OUT, I2 => G_5184GAT_OUT, O 
                           => G_5251GAT_OUT);
   G_5250GAT : Nor_gate port map( I1 => G_5184GAT_OUT, I2 => G_675GAT_OUT, O =>
                           G_5250GAT_OUT);
   G_5249GAT : Nor_gate port map( I1 => G_5124GAT_OUT, I2 => G_5184GAT_OUT, O 
                           => G_5249GAT_OUT);
   G_5246GAT : Nor_gate port map( I1 => G_5009GAT_OUT, I2 => G_5180GAT_OUT, O 
                           => G_5246GAT_OUT);
   G_5245GAT : Nor_gate port map( I1 => G_5180GAT_OUT, I2 => G_627GAT_OUT, O =>
                           G_5245GAT_OUT);
   G_5244GAT : Nor_gate port map( I1 => G_5121GAT_OUT, I2 => G_5180GAT_OUT, O 
                           => G_5244GAT_OUT);
   G_5241GAT : Nor_gate port map( I1 => G_5005GAT_OUT, I2 => G_5176GAT_OUT, O 
                           => G_5241GAT_OUT);
   G_5240GAT : Nor_gate port map( I1 => G_5176GAT_OUT, I2 => G_579GAT_OUT, O =>
                           G_5240GAT_OUT);
   G_5239GAT : Nor_gate port map( I1 => G_5118GAT_OUT, I2 => G_5176GAT_OUT, O 
                           => G_5239GAT_OUT);
   G_5236GAT : Nor_gate port map( I1 => G_5001GAT_OUT, I2 => G_5172GAT_OUT, O 
                           => G_5236GAT_OUT);
   G_5235GAT : Nor_gate port map( I1 => G_5172GAT_OUT, I2 => G_1257GAT_OUT, O 
                           => G_5235GAT_OUT);
   G_5234GAT : Nor_gate port map( I1 => G_5115GAT_OUT, I2 => G_5172GAT_OUT, O 
                           => G_5234GAT_OUT);
   G_5230GAT : Nor_gate port map( I1 => G_5169GAT_OUT, I2 => G_1209GAT_OUT, O 
                           => G_5230GAT_OUT);
   G_5227GAT : Nor_gate port map( I1 => G_5167GAT_OUT, I2 => G_5168GAT_OUT, O 
                           => G_5227GAT_OUT);
   G_5226GAT : Nor_gate port map( I1 => G_5163GAT_OUT, I2 => G_5103GAT_OUT, O 
                           => G_5226GAT_OUT);
   G_5225GAT : Nor_gate port map( I1 => G_5106GAT_OUT, I2 => G_5163GAT_OUT, O 
                           => G_5225GAT_OUT);
   G_5221GAT : Nor_gate port map( I1 => G_5160GAT_OUT, I2 => G_5157GAT_OUT, O 
                           => G_5221GAT_OUT);
   G_5218GAT : Nor_gate port map( I1 => G_5155GAT_OUT, I2 => G_5156GAT_OUT, O 
                           => G_5218GAT_OUT);
   G_5215GAT : Nor_gate port map( I1 => G_4980GAT_OUT, I2 => G_5151GAT_OUT, O 
                           => G_5215GAT_OUT);
   G_5214GAT : Nor_gate port map( I1 => G_5151GAT_OUT, I2 => G_1014GAT_OUT, O 
                           => G_5214GAT_OUT);
   G_5213GAT : Nor_gate port map( I1 => G_5094GAT_OUT, I2 => G_5151GAT_OUT, O 
                           => G_5213GAT_OUT);
   G_5209GAT : Nor_gate port map( I1 => G_5148GAT_OUT, I2 => G_966GAT_OUT, O =>
                           G_5209GAT_OUT);
   G_5206GAT : Nor_gate port map( I1 => G_5146GAT_OUT, I2 => G_5147GAT_OUT, O 
                           => G_5206GAT_OUT);
   G_5205GAT : Nor_gate port map( I1 => G_5142GAT_OUT, I2 => G_5082GAT_OUT, O 
                           => G_5205GAT_OUT);
   G_5204GAT : Nor_gate port map( I1 => G_5085GAT_OUT, I2 => G_5142GAT_OUT, O 
                           => G_5204GAT_OUT);
   G_5200GAT : Nor_gate port map( I1 => G_5139GAT_OUT, I2 => G_5136GAT_OUT, O 
                           => G_5200GAT_OUT);
   G_5197GAT : Nor_gate port map( I1 => G_5134GAT_OUT, I2 => G_5135GAT_OUT, O 
                           => G_5197GAT_OUT);
   G_5194GAT : Nor_gate port map( I1 => G_4959GAT_OUT, I2 => G_5130GAT_OUT, O 
                           => G_5194GAT_OUT);
   G_5193GAT : Nor_gate port map( I1 => G_5130GAT_OUT, I2 => G_771GAT_OUT, O =>
                           G_5193GAT_OUT);
   G_5192GAT : Nor_gate port map( I1 => G_5073GAT_OUT, I2 => G_5130GAT_OUT, O 
                           => G_5192GAT_OUT);
   G_5188GAT : Nor_gate port map( I1 => G_5127GAT_OUT, I2 => G_723GAT_OUT, O =>
                           G_5188GAT_OUT);
   G_5184GAT : Nor_gate port map( I1 => G_5124GAT_OUT, I2 => G_675GAT_OUT, O =>
                           G_5184GAT_OUT);
   G_5180GAT : Nor_gate port map( I1 => G_5121GAT_OUT, I2 => G_627GAT_OUT, O =>
                           G_5180GAT_OUT);
   G_5176GAT : Nor_gate port map( I1 => G_5118GAT_OUT, I2 => G_579GAT_OUT, O =>
                           G_5176GAT_OUT);
   G_5172GAT : Nor_gate port map( I1 => G_5115GAT_OUT, I2 => G_1257GAT_OUT, O 
                           => G_5172GAT_OUT);
   G_5169GAT : Nor_gate port map( I1 => G_5113GAT_OUT, I2 => G_5114GAT_OUT, O 
                           => G_5169GAT_OUT);
   G_5168GAT : Nor_gate port map( I1 => G_5109GAT_OUT, I2 => G_5053GAT_OUT, O 
                           => G_5168GAT_OUT);
   G_5167GAT : Nor_gate port map( I1 => G_5056GAT_OUT, I2 => G_5109GAT_OUT, O 
                           => G_5167GAT_OUT);
   G_5163GAT : Nor_gate port map( I1 => G_5106GAT_OUT, I2 => G_5103GAT_OUT, O 
                           => G_5163GAT_OUT);
   G_5160GAT : Nor_gate port map( I1 => G_5101GAT_OUT, I2 => G_5102GAT_OUT, O 
                           => G_5160GAT_OUT);
   G_5157GAT : Nor_gate port map( I1 => G_4928GAT_OUT, I2 => G_5097GAT_OUT, O 
                           => G_5157GAT_OUT);
   G_5156GAT : Nor_gate port map( I1 => G_5097GAT_OUT, I2 => G_1062GAT_OUT, O 
                           => G_5156GAT_OUT);
   G_5155GAT : Nor_gate port map( I1 => G_5044GAT_OUT, I2 => G_5097GAT_OUT, O 
                           => G_5155GAT_OUT);
   G_5151GAT : Nor_gate port map( I1 => G_5094GAT_OUT, I2 => G_1014GAT_OUT, O 
                           => G_5151GAT_OUT);
   G_5148GAT : Nor_gate port map( I1 => G_5092GAT_OUT, I2 => G_5093GAT_OUT, O 
                           => G_5148GAT_OUT);
   G_5147GAT : Nor_gate port map( I1 => G_5088GAT_OUT, I2 => G_5032GAT_OUT, O 
                           => G_5147GAT_OUT);
   G_5146GAT : Nor_gate port map( I1 => G_5035GAT_OUT, I2 => G_5088GAT_OUT, O 
                           => G_5146GAT_OUT);
   G_5142GAT : Nor_gate port map( I1 => G_5085GAT_OUT, I2 => G_5082GAT_OUT, O 
                           => G_5142GAT_OUT);
   G_5139GAT : Nor_gate port map( I1 => G_5080GAT_OUT, I2 => G_5081GAT_OUT, O 
                           => G_5139GAT_OUT);
   G_5136GAT : Nor_gate port map( I1 => G_4907GAT_OUT, I2 => G_5076GAT_OUT, O 
                           => G_5136GAT_OUT);
   G_5135GAT : Nor_gate port map( I1 => G_5076GAT_OUT, I2 => G_819GAT_OUT, O =>
                           G_5135GAT_OUT);
   G_5134GAT : Nor_gate port map( I1 => G_5023GAT_OUT, I2 => G_5076GAT_OUT, O 
                           => G_5134GAT_OUT);
   G_5130GAT : Nor_gate port map( I1 => G_5073GAT_OUT, I2 => G_771GAT_OUT, O =>
                           G_5130GAT_OUT);
   G_5127GAT : Nor_gate port map( I1 => G_5071GAT_OUT, I2 => G_5072GAT_OUT, O 
                           => G_5127GAT_OUT);
   G_5124GAT : Nor_gate port map( I1 => G_5069GAT_OUT, I2 => G_5070GAT_OUT, O 
                           => G_5124GAT_OUT);
   G_5121GAT : Nor_gate port map( I1 => G_5067GAT_OUT, I2 => G_5068GAT_OUT, O 
                           => G_5121GAT_OUT);
   G_5118GAT : Nor_gate port map( I1 => G_5065GAT_OUT, I2 => G_5066GAT_OUT, O 
                           => G_5118GAT_OUT);
   G_5115GAT : Nor_gate port map( I1 => G_5063GAT_OUT, I2 => G_5064GAT_OUT, O 
                           => G_5115GAT_OUT);
   G_5114GAT : Nor_gate port map( I1 => G_5059GAT_OUT, I2 => G_4995GAT_OUT, O 
                           => G_5114GAT_OUT);
   G_5113GAT : Nor_gate port map( I1 => G_4998GAT_OUT, I2 => G_5059GAT_OUT, O 
                           => G_5113GAT_OUT);
   G_5109GAT : Nor_gate port map( I1 => G_5056GAT_OUT, I2 => G_5053GAT_OUT, O 
                           => G_5109GAT_OUT);
   G_5106GAT : Nor_gate port map( I1 => G_5051GAT_OUT, I2 => G_5052GAT_OUT, O 
                           => G_5106GAT_OUT);
   G_5103GAT : Nor_gate port map( I1 => G_4866GAT_OUT, I2 => G_5047GAT_OUT, O 
                           => G_5103GAT_OUT);
   G_5102GAT : Nor_gate port map( I1 => G_5047GAT_OUT, I2 => G_1110GAT_OUT, O 
                           => G_5102GAT_OUT);
   G_5101GAT : Nor_gate port map( I1 => G_4986GAT_OUT, I2 => G_5047GAT_OUT, O 
                           => G_5101GAT_OUT);
   G_5097GAT : Nor_gate port map( I1 => G_5044GAT_OUT, I2 => G_1062GAT_OUT, O 
                           => G_5097GAT_OUT);
   G_5094GAT : Nor_gate port map( I1 => G_5042GAT_OUT, I2 => G_5043GAT_OUT, O 
                           => G_5094GAT_OUT);
   G_5093GAT : Nor_gate port map( I1 => G_5038GAT_OUT, I2 => G_4974GAT_OUT, O 
                           => G_5093GAT_OUT);
   G_5092GAT : Nor_gate port map( I1 => G_4977GAT_OUT, I2 => G_5038GAT_OUT, O 
                           => G_5092GAT_OUT);
   G_5088GAT : Nor_gate port map( I1 => G_5035GAT_OUT, I2 => G_5032GAT_OUT, O 
                           => G_5088GAT_OUT);
   G_5085GAT : Nor_gate port map( I1 => G_5030GAT_OUT, I2 => G_5031GAT_OUT, O 
                           => G_5085GAT_OUT);
   G_5082GAT : Nor_gate port map( I1 => G_4845GAT_OUT, I2 => G_5026GAT_OUT, O 
                           => G_5082GAT_OUT);
   G_5081GAT : Nor_gate port map( I1 => G_5026GAT_OUT, I2 => G_867GAT_OUT, O =>
                           G_5081GAT_OUT);
   G_5080GAT : Nor_gate port map( I1 => G_4965GAT_OUT, I2 => G_5026GAT_OUT, O 
                           => G_5080GAT_OUT);
   G_5076GAT : Nor_gate port map( I1 => G_5023GAT_OUT, I2 => G_819GAT_OUT, O =>
                           G_5076GAT_OUT);
   G_5073GAT : Nor_gate port map( I1 => G_5021GAT_OUT, I2 => G_5022GAT_OUT, O 
                           => G_5073GAT_OUT);
   G_5072GAT : Nor_gate port map( I1 => G_5017GAT_OUT, I2 => G_4896GAT_OUT, O 
                           => G_5072GAT_OUT);
   G_5071GAT : Nor_gate port map( I1 => G_4956GAT_OUT, I2 => G_5017GAT_OUT, O 
                           => G_5071GAT_OUT);
   G_5070GAT : Nor_gate port map( I1 => G_5013GAT_OUT, I2 => G_4891GAT_OUT, O 
                           => G_5070GAT_OUT);
   G_5069GAT : Nor_gate port map( I1 => G_4953GAT_OUT, I2 => G_5013GAT_OUT, O 
                           => G_5069GAT_OUT);
   G_5068GAT : Nor_gate port map( I1 => G_5009GAT_OUT, I2 => G_4886GAT_OUT, O 
                           => G_5068GAT_OUT);
   G_5067GAT : Nor_gate port map( I1 => G_4950GAT_OUT, I2 => G_5009GAT_OUT, O 
                           => G_5067GAT_OUT);
   G_5066GAT : Nor_gate port map( I1 => G_5005GAT_OUT, I2 => G_4881GAT_OUT, O 
                           => G_5066GAT_OUT);
   G_5065GAT : Nor_gate port map( I1 => G_4947GAT_OUT, I2 => G_5005GAT_OUT, O 
                           => G_5065GAT_OUT);
   G_5064GAT : Nor_gate port map( I1 => G_5001GAT_OUT, I2 => G_4943GAT_OUT, O 
                           => G_5064GAT_OUT);
   G_5063GAT : Nor_gate port map( I1 => G_1302GAT_OUT, I2 => G_5001GAT_OUT, O 
                           => G_5063GAT_OUT);
   G_5059GAT : Nor_gate port map( I1 => G_4998GAT_OUT, I2 => G_4995GAT_OUT, O 
                           => G_5059GAT_OUT);
   G_5056GAT : Nor_gate port map( I1 => G_4993GAT_OUT, I2 => G_4994GAT_OUT, O 
                           => G_5056GAT_OUT);
   G_5053GAT : Nor_gate port map( I1 => G_4808GAT_OUT, I2 => G_4989GAT_OUT, O 
                           => G_5053GAT_OUT);
   G_5052GAT : Nor_gate port map( I1 => G_4989GAT_OUT, I2 => G_1158GAT_OUT, O 
                           => G_5052GAT_OUT);
   G_5051GAT : Nor_gate port map( I1 => G_4934GAT_OUT, I2 => G_4989GAT_OUT, O 
                           => G_5051GAT_OUT);
   G_5047GAT : Nor_gate port map( I1 => G_4986GAT_OUT, I2 => G_1110GAT_OUT, O 
                           => G_5047GAT_OUT);
   G_5044GAT : Nor_gate port map( I1 => G_4984GAT_OUT, I2 => G_4985GAT_OUT, O 
                           => G_5044GAT_OUT);
   G_5043GAT : Nor_gate port map( I1 => G_4980GAT_OUT, I2 => G_4922GAT_OUT, O 
                           => G_5043GAT_OUT);
   G_5042GAT : Nor_gate port map( I1 => G_4925GAT_OUT, I2 => G_4980GAT_OUT, O 
                           => G_5042GAT_OUT);
   G_5038GAT : Nor_gate port map( I1 => G_4977GAT_OUT, I2 => G_4974GAT_OUT, O 
                           => G_5038GAT_OUT);
   G_5035GAT : Nor_gate port map( I1 => G_4972GAT_OUT, I2 => G_4973GAT_OUT, O 
                           => G_5035GAT_OUT);
   G_5032GAT : Nor_gate port map( I1 => G_4787GAT_OUT, I2 => G_4968GAT_OUT, O 
                           => G_5032GAT_OUT);
   G_5031GAT : Nor_gate port map( I1 => G_4968GAT_OUT, I2 => G_915GAT_OUT, O =>
                           G_5031GAT_OUT);
   G_5030GAT : Nor_gate port map( I1 => G_4913GAT_OUT, I2 => G_4968GAT_OUT, O 
                           => G_5030GAT_OUT);
   G_5026GAT : Nor_gate port map( I1 => G_4965GAT_OUT, I2 => G_867GAT_OUT, O =>
                           G_5026GAT_OUT);
   G_5023GAT : Nor_gate port map( I1 => G_4963GAT_OUT, I2 => G_4964GAT_OUT, O 
                           => G_5023GAT_OUT);
   G_5022GAT : Nor_gate port map( I1 => G_4959GAT_OUT, I2 => G_4901GAT_OUT, O 
                           => G_5022GAT_OUT);
   G_5021GAT : Nor_gate port map( I1 => G_4904GAT_OUT, I2 => G_4959GAT_OUT, O 
                           => G_5021GAT_OUT);
   G_5017GAT : Nor_gate port map( I1 => G_4956GAT_OUT, I2 => G_4896GAT_OUT, O 
                           => G_5017GAT_OUT);
   G_5013GAT : Nor_gate port map( I1 => G_4953GAT_OUT, I2 => G_4891GAT_OUT, O 
                           => G_5013GAT_OUT);
   G_5009GAT : Nor_gate port map( I1 => G_4950GAT_OUT, I2 => G_4886GAT_OUT, O 
                           => G_5009GAT_OUT);
   G_5005GAT : Nor_gate port map( I1 => G_4947GAT_OUT, I2 => G_4881GAT_OUT, O 
                           => G_5005GAT_OUT);
   G_5001GAT : Nor_gate port map( I1 => G_1302GAT_OUT, I2 => G_4943GAT_OUT, O 
                           => G_5001GAT_OUT);
   G_4998GAT : Nor_gate port map( I1 => G_4941GAT_OUT, I2 => G_4942GAT_OUT, O 
                           => G_4998GAT_OUT);
   G_4995GAT : Nor_gate port map( I1 => G_4754GAT_OUT, I2 => G_4937GAT_OUT, O 
                           => G_4995GAT_OUT);
   G_4994GAT : Nor_gate port map( I1 => G_4937GAT_OUT, I2 => G_1206GAT_OUT, O 
                           => G_4994GAT_OUT);
   G_4993GAT : Nor_gate port map( I1 => G_4872GAT_OUT, I2 => G_4937GAT_OUT, O 
                           => G_4993GAT_OUT);
   G_4989GAT : Nor_gate port map( I1 => G_4934GAT_OUT, I2 => G_1158GAT_OUT, O 
                           => G_4989GAT_OUT);
   G_4986GAT : Nor_gate port map( I1 => G_4932GAT_OUT, I2 => G_4933GAT_OUT, O 
                           => G_4986GAT_OUT);
   G_4985GAT : Nor_gate port map( I1 => G_4928GAT_OUT, I2 => G_4860GAT_OUT, O 
                           => G_4985GAT_OUT);
   G_4984GAT : Nor_gate port map( I1 => G_4863GAT_OUT, I2 => G_4928GAT_OUT, O 
                           => G_4984GAT_OUT);
   G_4980GAT : Nor_gate port map( I1 => G_4925GAT_OUT, I2 => G_4922GAT_OUT, O 
                           => G_4980GAT_OUT);
   G_4977GAT : Nor_gate port map( I1 => G_4920GAT_OUT, I2 => G_4921GAT_OUT, O 
                           => G_4977GAT_OUT);
   G_4974GAT : Nor_gate port map( I1 => G_4733GAT_OUT, I2 => G_4916GAT_OUT, O 
                           => G_4974GAT_OUT);
   G_4973GAT : Nor_gate port map( I1 => G_4916GAT_OUT, I2 => G_963GAT_OUT, O =>
                           G_4973GAT_OUT);
   G_4972GAT : Nor_gate port map( I1 => G_4851GAT_OUT, I2 => G_4916GAT_OUT, O 
                           => G_4972GAT_OUT);
   G_4968GAT : Nor_gate port map( I1 => G_4913GAT_OUT, I2 => G_915GAT_OUT, O =>
                           G_4968GAT_OUT);
   G_4965GAT : Nor_gate port map( I1 => G_4911GAT_OUT, I2 => G_4912GAT_OUT, O 
                           => G_4965GAT_OUT);
   G_4964GAT : Nor_gate port map( I1 => G_4907GAT_OUT, I2 => G_4839GAT_OUT, O 
                           => G_4964GAT_OUT);
   G_4963GAT : Nor_gate port map( I1 => G_4842GAT_OUT, I2 => G_4907GAT_OUT, O 
                           => G_4963GAT_OUT);
   G_4959GAT : Nor_gate port map( I1 => G_4904GAT_OUT, I2 => G_4901GAT_OUT, O 
                           => G_4959GAT_OUT);
   G_4956GAT : Nor_gate port map( I1 => G_4899GAT_OUT, I2 => G_4900GAT_OUT, O 
                           => G_4956GAT_OUT);
   G_4953GAT : Nor_gate port map( I1 => G_4894GAT_OUT, I2 => G_4895GAT_OUT, O 
                           => G_4953GAT_OUT);
   G_4950GAT : Nor_gate port map( I1 => G_4889GAT_OUT, I2 => G_4890GAT_OUT, O 
                           => G_4950GAT_OUT);
   G_4947GAT : Nor_gate port map( I1 => G_4884GAT_OUT, I2 => G_4885GAT_OUT, O 
                           => G_4947GAT_OUT);
   G_4943GAT : Nor_gate port map( I1 => G_4704GAT_OUT, I2 => G_4875GAT_OUT, O 
                           => G_4943GAT_OUT);
   G_4942GAT : Nor_gate port map( I1 => G_4875GAT_OUT, I2 => G_1254GAT_OUT, O 
                           => G_4942GAT_OUT);
   G_4941GAT : Nor_gate port map( I1 => G_4814GAT_OUT, I2 => G_4875GAT_OUT, O 
                           => G_4941GAT_OUT);
   G_4937GAT : Nor_gate port map( I1 => G_4872GAT_OUT, I2 => G_1206GAT_OUT, O 
                           => G_4937GAT_OUT);
   G_4934GAT : Nor_gate port map( I1 => G_4870GAT_OUT, I2 => G_4871GAT_OUT, O 
                           => G_4934GAT_OUT);
   G_4933GAT : Nor_gate port map( I1 => G_4866GAT_OUT, I2 => G_4802GAT_OUT, O 
                           => G_4933GAT_OUT);
   G_4932GAT : Nor_gate port map( I1 => G_4805GAT_OUT, I2 => G_4866GAT_OUT, O 
                           => G_4932GAT_OUT);
   G_4928GAT : Nor_gate port map( I1 => G_4863GAT_OUT, I2 => G_4860GAT_OUT, O 
                           => G_4928GAT_OUT);
   G_4925GAT : Nor_gate port map( I1 => G_4858GAT_OUT, I2 => G_4859GAT_OUT, O 
                           => G_4925GAT_OUT);
   G_4922GAT : Nor_gate port map( I1 => G_4683GAT_OUT, I2 => G_4854GAT_OUT, O 
                           => G_4922GAT_OUT);
   G_4921GAT : Nor_gate port map( I1 => G_4854GAT_OUT, I2 => G_1011GAT_OUT, O 
                           => G_4921GAT_OUT);
   G_4920GAT : Nor_gate port map( I1 => G_4793GAT_OUT, I2 => G_4854GAT_OUT, O 
                           => G_4920GAT_OUT);
   G_4916GAT : Nor_gate port map( I1 => G_4851GAT_OUT, I2 => G_963GAT_OUT, O =>
                           G_4916GAT_OUT);
   G_4913GAT : Nor_gate port map( I1 => G_4849GAT_OUT, I2 => G_4850GAT_OUT, O 
                           => G_4913GAT_OUT);
   G_4912GAT : Nor_gate port map( I1 => G_4845GAT_OUT, I2 => G_4781GAT_OUT, O 
                           => G_4912GAT_OUT);
   G_4911GAT : Nor_gate port map( I1 => G_4784GAT_OUT, I2 => G_4845GAT_OUT, O 
                           => G_4911GAT_OUT);
   G_4907GAT : Nor_gate port map( I1 => G_4842GAT_OUT, I2 => G_4839GAT_OUT, O 
                           => G_4907GAT_OUT);
   G_4904GAT : Nor_gate port map( I1 => G_4837GAT_OUT, I2 => G_4838GAT_OUT, O 
                           => G_4904GAT_OUT);
   G_4901GAT : Nor_gate port map( I1 => G_4662GAT_OUT, I2 => G_4833GAT_OUT, O 
                           => G_4901GAT_OUT);
   G_4900GAT : Nor_gate port map( I1 => G_4833GAT_OUT, I2 => G_768GAT_OUT, O =>
                           G_4900GAT_OUT);
   G_4899GAT : Nor_gate port map( I1 => G_4772GAT_OUT, I2 => G_4833GAT_OUT, O 
                           => G_4899GAT_OUT);
   G_4896GAT : Nor_gate port map( I1 => G_4658GAT_OUT, I2 => G_4829GAT_OUT, O 
                           => G_4896GAT_OUT);
   G_4895GAT : Nor_gate port map( I1 => G_4829GAT_OUT, I2 => G_720GAT_OUT, O =>
                           G_4895GAT_OUT);
   G_4894GAT : Nor_gate port map( I1 => G_4769GAT_OUT, I2 => G_4829GAT_OUT, O 
                           => G_4894GAT_OUT);
   G_4891GAT : Nor_gate port map( I1 => G_4654GAT_OUT, I2 => G_4825GAT_OUT, O 
                           => G_4891GAT_OUT);
   G_4890GAT : Nor_gate port map( I1 => G_4825GAT_OUT, I2 => G_672GAT_OUT, O =>
                           G_4890GAT_OUT);
   G_4889GAT : Nor_gate port map( I1 => G_4766GAT_OUT, I2 => G_4825GAT_OUT, O 
                           => G_4889GAT_OUT);
   G_4886GAT : Nor_gate port map( I1 => G_4650GAT_OUT, I2 => G_4821GAT_OUT, O 
                           => G_4886GAT_OUT);
   G_4885GAT : Nor_gate port map( I1 => G_4821GAT_OUT, I2 => G_624GAT_OUT, O =>
                           G_4885GAT_OUT);
   G_4884GAT : Nor_gate port map( I1 => G_4763GAT_OUT, I2 => G_4821GAT_OUT, O 
                           => G_4884GAT_OUT);
   G_4881GAT : Nor_gate port map( I1 => G_4646GAT_OUT, I2 => G_4817GAT_OUT, O 
                           => G_4881GAT_OUT);
   G_4880GAT : Nor_gate port map( I1 => G_4817GAT_OUT, I2 => G_576GAT_OUT, O =>
                           G_4880GAT_OUT);
   G_4879GAT : Nor_gate port map( I1 => G_4760GAT_OUT, I2 => G_4817GAT_OUT, O 
                           => G_4879GAT_OUT);
   G_4875GAT : Nor_gate port map( I1 => G_4814GAT_OUT, I2 => G_1254GAT_OUT, O 
                           => G_4875GAT_OUT);
   G_4872GAT : Nor_gate port map( I1 => G_4812GAT_OUT, I2 => G_4813GAT_OUT, O 
                           => G_4872GAT_OUT);
   G_4871GAT : Nor_gate port map( I1 => G_4808GAT_OUT, I2 => G_4748GAT_OUT, O 
                           => G_4871GAT_OUT);
   G_4870GAT : Nor_gate port map( I1 => G_4751GAT_OUT, I2 => G_4808GAT_OUT, O 
                           => G_4870GAT_OUT);
   G_4866GAT : Nor_gate port map( I1 => G_4805GAT_OUT, I2 => G_4802GAT_OUT, O 
                           => G_4866GAT_OUT);
   G_4863GAT : Nor_gate port map( I1 => G_4800GAT_OUT, I2 => G_4801GAT_OUT, O 
                           => G_4863GAT_OUT);
   G_4860GAT : Nor_gate port map( I1 => G_4628GAT_OUT, I2 => G_4796GAT_OUT, O 
                           => G_4860GAT_OUT);
   G_4859GAT : Nor_gate port map( I1 => G_4796GAT_OUT, I2 => G_1059GAT_OUT, O 
                           => G_4859GAT_OUT);
   G_4858GAT : Nor_gate port map( I1 => G_4739GAT_OUT, I2 => G_4796GAT_OUT, O 
                           => G_4858GAT_OUT);
   G_4854GAT : Nor_gate port map( I1 => G_4793GAT_OUT, I2 => G_1011GAT_OUT, O 
                           => G_4854GAT_OUT);
   G_4851GAT : Nor_gate port map( I1 => G_4791GAT_OUT, I2 => G_4792GAT_OUT, O 
                           => G_4851GAT_OUT);
   G_4850GAT : Nor_gate port map( I1 => G_4787GAT_OUT, I2 => G_4727GAT_OUT, O 
                           => G_4850GAT_OUT);
   G_4849GAT : Nor_gate port map( I1 => G_4730GAT_OUT, I2 => G_4787GAT_OUT, O 
                           => G_4849GAT_OUT);
   G_4845GAT : Nor_gate port map( I1 => G_4784GAT_OUT, I2 => G_4781GAT_OUT, O 
                           => G_4845GAT_OUT);
   G_4842GAT : Nor_gate port map( I1 => G_4779GAT_OUT, I2 => G_4780GAT_OUT, O 
                           => G_4842GAT_OUT);
   G_4839GAT : Nor_gate port map( I1 => G_4607GAT_OUT, I2 => G_4775GAT_OUT, O 
                           => G_4839GAT_OUT);
   G_4838GAT : Nor_gate port map( I1 => G_4775GAT_OUT, I2 => G_816GAT_OUT, O =>
                           G_4838GAT_OUT);
   G_4837GAT : Nor_gate port map( I1 => G_4718GAT_OUT, I2 => G_4775GAT_OUT, O 
                           => G_4837GAT_OUT);
   G_4833GAT : Nor_gate port map( I1 => G_4772GAT_OUT, I2 => G_768GAT_OUT, O =>
                           G_4833GAT_OUT);
   G_4829GAT : Nor_gate port map( I1 => G_4769GAT_OUT, I2 => G_720GAT_OUT, O =>
                           G_4829GAT_OUT);
   G_4825GAT : Nor_gate port map( I1 => G_4766GAT_OUT, I2 => G_672GAT_OUT, O =>
                           G_4825GAT_OUT);
   G_4821GAT : Nor_gate port map( I1 => G_4763GAT_OUT, I2 => G_624GAT_OUT, O =>
                           G_4821GAT_OUT);
   G_4817GAT : Nor_gate port map( I1 => G_4760GAT_OUT, I2 => G_576GAT_OUT, O =>
                           G_4817GAT_OUT);
   G_4814GAT : Nor_gate port map( I1 => G_4758GAT_OUT, I2 => G_4759GAT_OUT, O 
                           => G_4814GAT_OUT);
   G_4813GAT : Nor_gate port map( I1 => G_4754GAT_OUT, I2 => G_4698GAT_OUT, O 
                           => G_4813GAT_OUT);
   G_4812GAT : Nor_gate port map( I1 => G_4701GAT_OUT, I2 => G_4754GAT_OUT, O 
                           => G_4812GAT_OUT);
   G_4808GAT : Nor_gate port map( I1 => G_4751GAT_OUT, I2 => G_4748GAT_OUT, O 
                           => G_4808GAT_OUT);
   G_4805GAT : Nor_gate port map( I1 => G_4746GAT_OUT, I2 => G_4747GAT_OUT, O 
                           => G_4805GAT_OUT);
   G_4802GAT : Nor_gate port map( I1 => G_4578GAT_OUT, I2 => G_4742GAT_OUT, O 
                           => G_4802GAT_OUT);
   G_4801GAT : Nor_gate port map( I1 => G_4742GAT_OUT, I2 => G_1107GAT_OUT, O 
                           => G_4801GAT_OUT);
   G_4800GAT : Nor_gate port map( I1 => G_4689GAT_OUT, I2 => G_4742GAT_OUT, O 
                           => G_4800GAT_OUT);
   G_4796GAT : Nor_gate port map( I1 => G_4739GAT_OUT, I2 => G_1059GAT_OUT, O 
                           => G_4796GAT_OUT);
   G_4793GAT : Nor_gate port map( I1 => G_4737GAT_OUT, I2 => G_4738GAT_OUT, O 
                           => G_4793GAT_OUT);
   G_4792GAT : Nor_gate port map( I1 => G_4733GAT_OUT, I2 => G_4677GAT_OUT, O 
                           => G_4792GAT_OUT);
   G_4791GAT : Nor_gate port map( I1 => G_4680GAT_OUT, I2 => G_4733GAT_OUT, O 
                           => G_4791GAT_OUT);
   G_4787GAT : Nor_gate port map( I1 => G_4730GAT_OUT, I2 => G_4727GAT_OUT, O 
                           => G_4787GAT_OUT);
   G_4784GAT : Nor_gate port map( I1 => G_4725GAT_OUT, I2 => G_4726GAT_OUT, O 
                           => G_4784GAT_OUT);
   G_4781GAT : Nor_gate port map( I1 => G_4557GAT_OUT, I2 => G_4721GAT_OUT, O 
                           => G_4781GAT_OUT);
   G_4780GAT : Nor_gate port map( I1 => G_4721GAT_OUT, I2 => G_864GAT_OUT, O =>
                           G_4780GAT_OUT);
   G_4779GAT : Nor_gate port map( I1 => G_4668GAT_OUT, I2 => G_4721GAT_OUT, O 
                           => G_4779GAT_OUT);
   G_4775GAT : Nor_gate port map( I1 => G_4718GAT_OUT, I2 => G_816GAT_OUT, O =>
                           G_4775GAT_OUT);
   G_4772GAT : Nor_gate port map( I1 => G_4716GAT_OUT, I2 => G_4717GAT_OUT, O 
                           => G_4772GAT_OUT);
   G_4769GAT : Nor_gate port map( I1 => G_4714GAT_OUT, I2 => G_4715GAT_OUT, O 
                           => G_4769GAT_OUT);
   G_4766GAT : Nor_gate port map( I1 => G_4712GAT_OUT, I2 => G_4713GAT_OUT, O 
                           => G_4766GAT_OUT);
   G_4763GAT : Nor_gate port map( I1 => G_4710GAT_OUT, I2 => G_4711GAT_OUT, O 
                           => G_4763GAT_OUT);
   G_4760GAT : Nor_gate port map( I1 => G_4708GAT_OUT, I2 => G_4709GAT_OUT, O 
                           => G_4760GAT_OUT);
   G_4759GAT : Nor_gate port map( I1 => G_4704GAT_OUT, I2 => G_4643GAT_OUT, O 
                           => G_4759GAT_OUT);
   G_4758GAT : Nor_gate port map( I1 => G_1299GAT_OUT, I2 => G_4704GAT_OUT, O 
                           => G_4758GAT_OUT);
   G_4754GAT : Nor_gate port map( I1 => G_4701GAT_OUT, I2 => G_4698GAT_OUT, O 
                           => G_4754GAT_OUT);
   G_4751GAT : Nor_gate port map( I1 => G_4696GAT_OUT, I2 => G_4697GAT_OUT, O 
                           => G_4751GAT_OUT);
   G_4748GAT : Nor_gate port map( I1 => G_4515GAT_OUT, I2 => G_4692GAT_OUT, O 
                           => G_4748GAT_OUT);
   G_4747GAT : Nor_gate port map( I1 => G_4692GAT_OUT, I2 => G_1155GAT_OUT, O 
                           => G_4747GAT_OUT);
   G_4746GAT : Nor_gate port map( I1 => G_4634GAT_OUT, I2 => G_4692GAT_OUT, O 
                           => G_4746GAT_OUT);
   G_4742GAT : Nor_gate port map( I1 => G_4689GAT_OUT, I2 => G_1107GAT_OUT, O 
                           => G_4742GAT_OUT);
   G_4739GAT : Nor_gate port map( I1 => G_4687GAT_OUT, I2 => G_4688GAT_OUT, O 
                           => G_4739GAT_OUT);
   G_4738GAT : Nor_gate port map( I1 => G_4683GAT_OUT, I2 => G_4622GAT_OUT, O 
                           => G_4738GAT_OUT);
   G_4737GAT : Nor_gate port map( I1 => G_4625GAT_OUT, I2 => G_4683GAT_OUT, O 
                           => G_4737GAT_OUT);
   G_4733GAT : Nor_gate port map( I1 => G_4680GAT_OUT, I2 => G_4677GAT_OUT, O 
                           => G_4733GAT_OUT);
   G_4730GAT : Nor_gate port map( I1 => G_4675GAT_OUT, I2 => G_4676GAT_OUT, O 
                           => G_4730GAT_OUT);
   G_4727GAT : Nor_gate port map( I1 => G_4494GAT_OUT, I2 => G_4671GAT_OUT, O 
                           => G_4727GAT_OUT);
   G_4726GAT : Nor_gate port map( I1 => G_4671GAT_OUT, I2 => G_912GAT_OUT, O =>
                           G_4726GAT_OUT);
   G_4725GAT : Nor_gate port map( I1 => G_4613GAT_OUT, I2 => G_4671GAT_OUT, O 
                           => G_4725GAT_OUT);
   G_4721GAT : Nor_gate port map( I1 => G_4668GAT_OUT, I2 => G_864GAT_OUT, O =>
                           G_4721GAT_OUT);
   G_4718GAT : Nor_gate port map( I1 => G_4666GAT_OUT, I2 => G_4667GAT_OUT, O 
                           => G_4718GAT_OUT);
   G_4717GAT : Nor_gate port map( I1 => G_4662GAT_OUT, I2 => G_4546GAT_OUT, O 
                           => G_4717GAT_OUT);
   G_4716GAT : Nor_gate port map( I1 => G_4604GAT_OUT, I2 => G_4662GAT_OUT, O 
                           => G_4716GAT_OUT);
   G_4715GAT : Nor_gate port map( I1 => G_4658GAT_OUT, I2 => G_4541GAT_OUT, O 
                           => G_4715GAT_OUT);
   G_4714GAT : Nor_gate port map( I1 => G_4601GAT_OUT, I2 => G_4658GAT_OUT, O 
                           => G_4714GAT_OUT);
   G_4713GAT : Nor_gate port map( I1 => G_4654GAT_OUT, I2 => G_4536GAT_OUT, O 
                           => G_4713GAT_OUT);
   G_4712GAT : Nor_gate port map( I1 => G_4598GAT_OUT, I2 => G_4654GAT_OUT, O 
                           => G_4712GAT_OUT);
   G_4711GAT : Nor_gate port map( I1 => G_4650GAT_OUT, I2 => G_4531GAT_OUT, O 
                           => G_4711GAT_OUT);
   G_4710GAT : Nor_gate port map( I1 => G_4595GAT_OUT, I2 => G_4650GAT_OUT, O 
                           => G_4710GAT_OUT);
   G_4709GAT : Nor_gate port map( I1 => G_4646GAT_OUT, I2 => G_4526GAT_OUT, O 
                           => G_4709GAT_OUT);
   G_4708GAT : Nor_gate port map( I1 => G_4592GAT_OUT, I2 => G_4646GAT_OUT, O 
                           => G_4708GAT_OUT);
   G_4704GAT : Nor_gate port map( I1 => G_1299GAT_OUT, I2 => G_4643GAT_OUT, O 
                           => G_4704GAT_OUT);
   G_4701GAT : Nor_gate port map( I1 => G_4641GAT_OUT, I2 => G_4642GAT_OUT, O 
                           => G_4701GAT_OUT);
   G_4698GAT : Nor_gate port map( I1 => G_4456GAT_OUT, I2 => G_4637GAT_OUT, O 
                           => G_4698GAT_OUT);
   G_4697GAT : Nor_gate port map( I1 => G_4637GAT_OUT, I2 => G_1203GAT_OUT, O 
                           => G_4697GAT_OUT);
   G_4696GAT : Nor_gate port map( I1 => G_4584GAT_OUT, I2 => G_4637GAT_OUT, O 
                           => G_4696GAT_OUT);
   G_4692GAT : Nor_gate port map( I1 => G_4634GAT_OUT, I2 => G_1155GAT_OUT, O 
                           => G_4692GAT_OUT);
   G_4689GAT : Nor_gate port map( I1 => G_4632GAT_OUT, I2 => G_4633GAT_OUT, O 
                           => G_4689GAT_OUT);
   G_4688GAT : Nor_gate port map( I1 => G_4628GAT_OUT, I2 => G_4572GAT_OUT, O 
                           => G_4688GAT_OUT);
   G_4687GAT : Nor_gate port map( I1 => G_4575GAT_OUT, I2 => G_4628GAT_OUT, O 
                           => G_4687GAT_OUT);
   G_4683GAT : Nor_gate port map( I1 => G_4625GAT_OUT, I2 => G_4622GAT_OUT, O 
                           => G_4683GAT_OUT);
   G_4680GAT : Nor_gate port map( I1 => G_4620GAT_OUT, I2 => G_4621GAT_OUT, O 
                           => G_4680GAT_OUT);
   G_4677GAT : Nor_gate port map( I1 => G_4435GAT_OUT, I2 => G_4616GAT_OUT, O 
                           => G_4677GAT_OUT);
   G_4676GAT : Nor_gate port map( I1 => G_4616GAT_OUT, I2 => G_960GAT_OUT, O =>
                           G_4676GAT_OUT);
   G_4675GAT : Nor_gate port map( I1 => G_4563GAT_OUT, I2 => G_4616GAT_OUT, O 
                           => G_4675GAT_OUT);
   G_4671GAT : Nor_gate port map( I1 => G_4613GAT_OUT, I2 => G_912GAT_OUT, O =>
                           G_4671GAT_OUT);
   G_4668GAT : Nor_gate port map( I1 => G_4611GAT_OUT, I2 => G_4612GAT_OUT, O 
                           => G_4668GAT_OUT);
   G_4667GAT : Nor_gate port map( I1 => G_4607GAT_OUT, I2 => G_4551GAT_OUT, O 
                           => G_4667GAT_OUT);
   G_4666GAT : Nor_gate port map( I1 => G_4554GAT_OUT, I2 => G_4607GAT_OUT, O 
                           => G_4666GAT_OUT);
   G_4662GAT : Nor_gate port map( I1 => G_4604GAT_OUT, I2 => G_4546GAT_OUT, O 
                           => G_4662GAT_OUT);
   G_4658GAT : Nor_gate port map( I1 => G_4601GAT_OUT, I2 => G_4541GAT_OUT, O 
                           => G_4658GAT_OUT);
   G_4654GAT : Nor_gate port map( I1 => G_4598GAT_OUT, I2 => G_4536GAT_OUT, O 
                           => G_4654GAT_OUT);
   G_4650GAT : Nor_gate port map( I1 => G_4595GAT_OUT, I2 => G_4531GAT_OUT, O 
                           => G_4650GAT_OUT);
   G_4646GAT : Nor_gate port map( I1 => G_4592GAT_OUT, I2 => G_4526GAT_OUT, O 
                           => G_4646GAT_OUT);
   G_4643GAT : Nor_gate port map( I1 => G_4401GAT_OUT, I2 => G_4587GAT_OUT, O 
                           => G_4643GAT_OUT);
   G_4642GAT : Nor_gate port map( I1 => G_4587GAT_OUT, I2 => G_1251GAT_OUT, O 
                           => G_4642GAT_OUT);
   G_4641GAT : Nor_gate port map( I1 => G_4521GAT_OUT, I2 => G_4587GAT_OUT, O 
                           => G_4641GAT_OUT);
   G_4637GAT : Nor_gate port map( I1 => G_4584GAT_OUT, I2 => G_1203GAT_OUT, O 
                           => G_4637GAT_OUT);
   G_4634GAT : Nor_gate port map( I1 => G_4582GAT_OUT, I2 => G_4583GAT_OUT, O 
                           => G_4634GAT_OUT);
   G_4633GAT : Nor_gate port map( I1 => G_4578GAT_OUT, I2 => G_4509GAT_OUT, O 
                           => G_4633GAT_OUT);
   G_4632GAT : Nor_gate port map( I1 => G_4512GAT_OUT, I2 => G_4578GAT_OUT, O 
                           => G_4632GAT_OUT);
   G_4628GAT : Nor_gate port map( I1 => G_4575GAT_OUT, I2 => G_4572GAT_OUT, O 
                           => G_4628GAT_OUT);
   G_4625GAT : Nor_gate port map( I1 => G_4570GAT_OUT, I2 => G_4571GAT_OUT, O 
                           => G_4625GAT_OUT);
   G_4622GAT : Nor_gate port map( I1 => G_4380GAT_OUT, I2 => G_4566GAT_OUT, O 
                           => G_4622GAT_OUT);
   G_4621GAT : Nor_gate port map( I1 => G_4566GAT_OUT, I2 => G_1008GAT_OUT, O 
                           => G_4621GAT_OUT);
   G_4620GAT : Nor_gate port map( I1 => G_4500GAT_OUT, I2 => G_4566GAT_OUT, O 
                           => G_4620GAT_OUT);
   G_4616GAT : Nor_gate port map( I1 => G_4563GAT_OUT, I2 => G_960GAT_OUT, O =>
                           G_4616GAT_OUT);
   G_4613GAT : Nor_gate port map( I1 => G_4561GAT_OUT, I2 => G_4562GAT_OUT, O 
                           => G_4613GAT_OUT);
   G_4612GAT : Nor_gate port map( I1 => G_4557GAT_OUT, I2 => G_4488GAT_OUT, O 
                           => G_4612GAT_OUT);
   G_4611GAT : Nor_gate port map( I1 => G_4491GAT_OUT, I2 => G_4557GAT_OUT, O 
                           => G_4611GAT_OUT);
   G_4607GAT : Nor_gate port map( I1 => G_4554GAT_OUT, I2 => G_4551GAT_OUT, O 
                           => G_4607GAT_OUT);
   G_4604GAT : Nor_gate port map( I1 => G_4549GAT_OUT, I2 => G_4550GAT_OUT, O 
                           => G_4604GAT_OUT);
   G_4601GAT : Nor_gate port map( I1 => G_4544GAT_OUT, I2 => G_4545GAT_OUT, O 
                           => G_4601GAT_OUT);
   G_4598GAT : Nor_gate port map( I1 => G_4539GAT_OUT, I2 => G_4540GAT_OUT, O 
                           => G_4598GAT_OUT);
   G_4595GAT : Nor_gate port map( I1 => G_4534GAT_OUT, I2 => G_4535GAT_OUT, O 
                           => G_4595GAT_OUT);
   G_4592GAT : Nor_gate port map( I1 => G_4529GAT_OUT, I2 => G_4530GAT_OUT, O 
                           => G_4592GAT_OUT);
   G_4587GAT : Nor_gate port map( I1 => G_4521GAT_OUT, I2 => G_1251GAT_OUT, O 
                           => G_4587GAT_OUT);
   G_4584GAT : Nor_gate port map( I1 => G_4519GAT_OUT, I2 => G_4520GAT_OUT, O 
                           => G_4584GAT_OUT);
   G_4583GAT : Nor_gate port map( I1 => G_4515GAT_OUT, I2 => G_4450GAT_OUT, O 
                           => G_4583GAT_OUT);
   G_4582GAT : Nor_gate port map( I1 => G_4453GAT_OUT, I2 => G_4515GAT_OUT, O 
                           => G_4582GAT_OUT);
   G_4578GAT : Nor_gate port map( I1 => G_4512GAT_OUT, I2 => G_4509GAT_OUT, O 
                           => G_4578GAT_OUT);
   G_4575GAT : Nor_gate port map( I1 => G_4507GAT_OUT, I2 => G_4508GAT_OUT, O 
                           => G_4575GAT_OUT);
   G_4572GAT : Nor_gate port map( I1 => G_4335GAT_OUT, I2 => G_4503GAT_OUT, O 
                           => G_4572GAT_OUT);
   G_4571GAT : Nor_gate port map( I1 => G_4503GAT_OUT, I2 => G_1056GAT_OUT, O 
                           => G_4571GAT_OUT);
   G_4570GAT : Nor_gate port map( I1 => G_4441GAT_OUT, I2 => G_4503GAT_OUT, O 
                           => G_4570GAT_OUT);
   G_4566GAT : Nor_gate port map( I1 => G_4500GAT_OUT, I2 => G_1008GAT_OUT, O 
                           => G_4566GAT_OUT);
   G_4563GAT : Nor_gate port map( I1 => G_4498GAT_OUT, I2 => G_4499GAT_OUT, O 
                           => G_4563GAT_OUT);
   G_4562GAT : Nor_gate port map( I1 => G_4494GAT_OUT, I2 => G_4429GAT_OUT, O 
                           => G_4562GAT_OUT);
   G_4561GAT : Nor_gate port map( I1 => G_4432GAT_OUT, I2 => G_4494GAT_OUT, O 
                           => G_4561GAT_OUT);
   G_4557GAT : Nor_gate port map( I1 => G_4491GAT_OUT, I2 => G_4488GAT_OUT, O 
                           => G_4557GAT_OUT);
   G_4554GAT : Nor_gate port map( I1 => G_4486GAT_OUT, I2 => G_4487GAT_OUT, O 
                           => G_4554GAT_OUT);
   G_4551GAT : Nor_gate port map( I1 => G_4314GAT_OUT, I2 => G_4482GAT_OUT, O 
                           => G_4551GAT_OUT);
   G_4550GAT : Nor_gate port map( I1 => G_4482GAT_OUT, I2 => G_813GAT_OUT, O =>
                           G_4550GAT_OUT);
   G_4549GAT : Nor_gate port map( I1 => G_4420GAT_OUT, I2 => G_4482GAT_OUT, O 
                           => G_4549GAT_OUT);
   G_4546GAT : Nor_gate port map( I1 => G_4310GAT_OUT, I2 => G_4478GAT_OUT, O 
                           => G_4546GAT_OUT);
   G_4545GAT : Nor_gate port map( I1 => G_4478GAT_OUT, I2 => G_765GAT_OUT, O =>
                           G_4545GAT_OUT);
   G_4544GAT : Nor_gate port map( I1 => G_4417GAT_OUT, I2 => G_4478GAT_OUT, O 
                           => G_4544GAT_OUT);
   G_4541GAT : Nor_gate port map( I1 => G_4306GAT_OUT, I2 => G_4474GAT_OUT, O 
                           => G_4541GAT_OUT);
   G_4540GAT : Nor_gate port map( I1 => G_4474GAT_OUT, I2 => G_717GAT_OUT, O =>
                           G_4540GAT_OUT);
   G_4539GAT : Nor_gate port map( I1 => G_4414GAT_OUT, I2 => G_4474GAT_OUT, O 
                           => G_4539GAT_OUT);
   G_4536GAT : Nor_gate port map( I1 => G_4302GAT_OUT, I2 => G_4470GAT_OUT, O 
                           => G_4536GAT_OUT);
   G_4535GAT : Nor_gate port map( I1 => G_4470GAT_OUT, I2 => G_669GAT_OUT, O =>
                           G_4535GAT_OUT);
   G_4534GAT : Nor_gate port map( I1 => G_4411GAT_OUT, I2 => G_4470GAT_OUT, O 
                           => G_4534GAT_OUT);
   G_4531GAT : Nor_gate port map( I1 => G_4298GAT_OUT, I2 => G_4466GAT_OUT, O 
                           => G_4531GAT_OUT);
   G_4530GAT : Nor_gate port map( I1 => G_4466GAT_OUT, I2 => G_621GAT_OUT, O =>
                           G_4530GAT_OUT);
   G_4529GAT : Nor_gate port map( I1 => G_4408GAT_OUT, I2 => G_4466GAT_OUT, O 
                           => G_4529GAT_OUT);
   G_4526GAT : Nor_gate port map( I1 => G_4294GAT_OUT, I2 => G_4462GAT_OUT, O 
                           => G_4526GAT_OUT);
   G_4525GAT : Nor_gate port map( I1 => G_4462GAT_OUT, I2 => G_573GAT_OUT, O =>
                           G_4525GAT_OUT);
   G_4524GAT : Nor_gate port map( I1 => G_4405GAT_OUT, I2 => G_4462GAT_OUT, O 
                           => G_4524GAT_OUT);
   G_4521GAT : Nor_gate port map( I1 => G_4460GAT_OUT, I2 => G_4461GAT_OUT, O 
                           => G_4521GAT_OUT);
   G_4520GAT : Nor_gate port map( I1 => G_4456GAT_OUT, I2 => G_4395GAT_OUT, O 
                           => G_4520GAT_OUT);
   G_4519GAT : Nor_gate port map( I1 => G_4398GAT_OUT, I2 => G_4456GAT_OUT, O 
                           => G_4519GAT_OUT);
   G_4515GAT : Nor_gate port map( I1 => G_4453GAT_OUT, I2 => G_4450GAT_OUT, O 
                           => G_4515GAT_OUT);
   G_4512GAT : Nor_gate port map( I1 => G_4448GAT_OUT, I2 => G_4449GAT_OUT, O 
                           => G_4512GAT_OUT);
   G_4509GAT : Nor_gate port map( I1 => G_4281GAT_OUT, I2 => G_4444GAT_OUT, O 
                           => G_4509GAT_OUT);
   G_4508GAT : Nor_gate port map( I1 => G_4444GAT_OUT, I2 => G_1104GAT_OUT, O 
                           => G_4508GAT_OUT);
   G_4507GAT : Nor_gate port map( I1 => G_4386GAT_OUT, I2 => G_4444GAT_OUT, O 
                           => G_4507GAT_OUT);
   G_4503GAT : Nor_gate port map( I1 => G_4441GAT_OUT, I2 => G_1056GAT_OUT, O 
                           => G_4503GAT_OUT);
   G_4500GAT : Nor_gate port map( I1 => G_4439GAT_OUT, I2 => G_4440GAT_OUT, O 
                           => G_4500GAT_OUT);
   G_4499GAT : Nor_gate port map( I1 => G_4435GAT_OUT, I2 => G_4374GAT_OUT, O 
                           => G_4499GAT_OUT);
   G_4498GAT : Nor_gate port map( I1 => G_4377GAT_OUT, I2 => G_4435GAT_OUT, O 
                           => G_4498GAT_OUT);
   G_4494GAT : Nor_gate port map( I1 => G_4432GAT_OUT, I2 => G_4429GAT_OUT, O 
                           => G_4494GAT_OUT);
   G_4491GAT : Nor_gate port map( I1 => G_4427GAT_OUT, I2 => G_4428GAT_OUT, O 
                           => G_4491GAT_OUT);
   G_4488GAT : Nor_gate port map( I1 => G_4260GAT_OUT, I2 => G_4423GAT_OUT, O 
                           => G_4488GAT_OUT);
   G_4487GAT : Nor_gate port map( I1 => G_4423GAT_OUT, I2 => G_861GAT_OUT, O =>
                           G_4487GAT_OUT);
   G_4486GAT : Nor_gate port map( I1 => G_4365GAT_OUT, I2 => G_4423GAT_OUT, O 
                           => G_4486GAT_OUT);
   G_4482GAT : Nor_gate port map( I1 => G_4420GAT_OUT, I2 => G_813GAT_OUT, O =>
                           G_4482GAT_OUT);
   G_4478GAT : Nor_gate port map( I1 => G_4417GAT_OUT, I2 => G_765GAT_OUT, O =>
                           G_4478GAT_OUT);
   G_4474GAT : Nor_gate port map( I1 => G_4414GAT_OUT, I2 => G_717GAT_OUT, O =>
                           G_4474GAT_OUT);
   G_4470GAT : Nor_gate port map( I1 => G_4411GAT_OUT, I2 => G_669GAT_OUT, O =>
                           G_4470GAT_OUT);
   G_4466GAT : Nor_gate port map( I1 => G_4408GAT_OUT, I2 => G_621GAT_OUT, O =>
                           G_4466GAT_OUT);
   G_4462GAT : Nor_gate port map( I1 => G_4405GAT_OUT, I2 => G_573GAT_OUT, O =>
                           G_4462GAT_OUT);
   G_4461GAT : Nor_gate port map( I1 => G_4401GAT_OUT, I2 => G_4350GAT_OUT, O 
                           => G_4461GAT_OUT);
   G_4460GAT : Nor_gate port map( I1 => G_1296GAT_OUT, I2 => G_4401GAT_OUT, O 
                           => G_4460GAT_OUT);
   G_4456GAT : Nor_gate port map( I1 => G_4398GAT_OUT, I2 => G_4395GAT_OUT, O 
                           => G_4456GAT_OUT);
   G_4453GAT : Nor_gate port map( I1 => G_4393GAT_OUT, I2 => G_4394GAT_OUT, O 
                           => G_4453GAT_OUT);
   G_4450GAT : Nor_gate port map( I1 => G_4232GAT_OUT, I2 => G_4389GAT_OUT, O 
                           => G_4450GAT_OUT);
   G_4449GAT : Nor_gate port map( I1 => G_4389GAT_OUT, I2 => G_1152GAT_OUT, O 
                           => G_4449GAT_OUT);
   G_4448GAT : Nor_gate port map( I1 => G_4341GAT_OUT, I2 => G_4389GAT_OUT, O 
                           => G_4448GAT_OUT);
   G_4444GAT : Nor_gate port map( I1 => G_4386GAT_OUT, I2 => G_1104GAT_OUT, O 
                           => G_4444GAT_OUT);
   G_4441GAT : Nor_gate port map( I1 => G_4384GAT_OUT, I2 => G_4385GAT_OUT, O 
                           => G_4441GAT_OUT);
   G_4440GAT : Nor_gate port map( I1 => G_4380GAT_OUT, I2 => G_4329GAT_OUT, O 
                           => G_4440GAT_OUT);
   G_4439GAT : Nor_gate port map( I1 => G_4332GAT_OUT, I2 => G_4380GAT_OUT, O 
                           => G_4439GAT_OUT);
   G_4435GAT : Nor_gate port map( I1 => G_4377GAT_OUT, I2 => G_4374GAT_OUT, O 
                           => G_4435GAT_OUT);
   G_4432GAT : Nor_gate port map( I1 => G_4372GAT_OUT, I2 => G_4373GAT_OUT, O 
                           => G_4432GAT_OUT);
   G_4429GAT : Nor_gate port map( I1 => G_4211GAT_OUT, I2 => G_4368GAT_OUT, O 
                           => G_4429GAT_OUT);
   G_4428GAT : Nor_gate port map( I1 => G_4368GAT_OUT, I2 => G_909GAT_OUT, O =>
                           G_4428GAT_OUT);
   G_4427GAT : Nor_gate port map( I1 => G_4320GAT_OUT, I2 => G_4368GAT_OUT, O 
                           => G_4427GAT_OUT);
   G_4423GAT : Nor_gate port map( I1 => G_4365GAT_OUT, I2 => G_861GAT_OUT, O =>
                           G_4423GAT_OUT);
   G_4420GAT : Nor_gate port map( I1 => G_4363GAT_OUT, I2 => G_4364GAT_OUT, O 
                           => G_4420GAT_OUT);
   G_4417GAT : Nor_gate port map( I1 => G_4361GAT_OUT, I2 => G_4362GAT_OUT, O 
                           => G_4417GAT_OUT);
   G_4414GAT : Nor_gate port map( I1 => G_4359GAT_OUT, I2 => G_4360GAT_OUT, O 
                           => G_4414GAT_OUT);
   G_4411GAT : Nor_gate port map( I1 => G_4357GAT_OUT, I2 => G_4358GAT_OUT, O 
                           => G_4411GAT_OUT);
   G_4408GAT : Nor_gate port map( I1 => G_4355GAT_OUT, I2 => G_4356GAT_OUT, O 
                           => G_4408GAT_OUT);
   G_4405GAT : Nor_gate port map( I1 => G_4353GAT_OUT, I2 => G_4354GAT_OUT, O 
                           => G_4405GAT_OUT);
   G_4401GAT : Nor_gate port map( I1 => G_1296GAT_OUT, I2 => G_4350GAT_OUT, O 
                           => G_4401GAT_OUT);
   G_4398GAT : Nor_gate port map( I1 => G_4348GAT_OUT, I2 => G_4349GAT_OUT, O 
                           => G_4398GAT_OUT);
   G_4395GAT : Nor_gate port map( I1 => G_4167GAT_OUT, I2 => G_4344GAT_OUT, O 
                           => G_4395GAT_OUT);
   G_4394GAT : Nor_gate port map( I1 => G_4344GAT_OUT, I2 => G_1200GAT_OUT, O 
                           => G_4394GAT_OUT);
   G_4393GAT : Nor_gate port map( I1 => G_4287GAT_OUT, I2 => G_4344GAT_OUT, O 
                           => G_4393GAT_OUT);
   G_4389GAT : Nor_gate port map( I1 => G_4341GAT_OUT, I2 => G_1152GAT_OUT, O 
                           => G_4389GAT_OUT);
   G_4386GAT : Nor_gate port map( I1 => G_4339GAT_OUT, I2 => G_4340GAT_OUT, O 
                           => G_4386GAT_OUT);
   G_4385GAT : Nor_gate port map( I1 => G_4335GAT_OUT, I2 => G_4275GAT_OUT, O 
                           => G_4385GAT_OUT);
   G_4384GAT : Nor_gate port map( I1 => G_4278GAT_OUT, I2 => G_4335GAT_OUT, O 
                           => G_4384GAT_OUT);
   G_4380GAT : Nor_gate port map( I1 => G_4332GAT_OUT, I2 => G_4329GAT_OUT, O 
                           => G_4380GAT_OUT);
   G_4377GAT : Nor_gate port map( I1 => G_4327GAT_OUT, I2 => G_4328GAT_OUT, O 
                           => G_4377GAT_OUT);
   G_4374GAT : Nor_gate port map( I1 => G_4146GAT_OUT, I2 => G_4323GAT_OUT, O 
                           => G_4374GAT_OUT);
   G_4373GAT : Nor_gate port map( I1 => G_4323GAT_OUT, I2 => G_957GAT_OUT, O =>
                           G_4373GAT_OUT);
   G_4372GAT : Nor_gate port map( I1 => G_4266GAT_OUT, I2 => G_4323GAT_OUT, O 
                           => G_4372GAT_OUT);
   G_4368GAT : Nor_gate port map( I1 => G_4320GAT_OUT, I2 => G_909GAT_OUT, O =>
                           G_4368GAT_OUT);
   G_4365GAT : Nor_gate port map( I1 => G_4318GAT_OUT, I2 => G_4319GAT_OUT, O 
                           => G_4365GAT_OUT);
   G_4364GAT : Nor_gate port map( I1 => G_4314GAT_OUT, I2 => G_4200GAT_OUT, O 
                           => G_4364GAT_OUT);
   G_4363GAT : Nor_gate port map( I1 => G_4257GAT_OUT, I2 => G_4314GAT_OUT, O 
                           => G_4363GAT_OUT);
   G_4362GAT : Nor_gate port map( I1 => G_4310GAT_OUT, I2 => G_4195GAT_OUT, O 
                           => G_4362GAT_OUT);
   G_4361GAT : Nor_gate port map( I1 => G_4254GAT_OUT, I2 => G_4310GAT_OUT, O 
                           => G_4361GAT_OUT);
   G_4360GAT : Nor_gate port map( I1 => G_4306GAT_OUT, I2 => G_4190GAT_OUT, O 
                           => G_4360GAT_OUT);
   G_4359GAT : Nor_gate port map( I1 => G_4251GAT_OUT, I2 => G_4306GAT_OUT, O 
                           => G_4359GAT_OUT);
   G_4358GAT : Nor_gate port map( I1 => G_4302GAT_OUT, I2 => G_4185GAT_OUT, O 
                           => G_4358GAT_OUT);
   G_4357GAT : Nor_gate port map( I1 => G_4248GAT_OUT, I2 => G_4302GAT_OUT, O 
                           => G_4357GAT_OUT);
   G_4356GAT : Nor_gate port map( I1 => G_4298GAT_OUT, I2 => G_4180GAT_OUT, O 
                           => G_4356GAT_OUT);
   G_4355GAT : Nor_gate port map( I1 => G_4245GAT_OUT, I2 => G_4298GAT_OUT, O 
                           => G_4355GAT_OUT);
   G_4354GAT : Nor_gate port map( I1 => G_4294GAT_OUT, I2 => G_4175GAT_OUT, O 
                           => G_4354GAT_OUT);
   G_4353GAT : Nor_gate port map( I1 => G_4242GAT_OUT, I2 => G_4294GAT_OUT, O 
                           => G_4353GAT_OUT);
   G_4350GAT : Nor_gate port map( I1 => G_4106GAT_OUT, I2 => G_4290GAT_OUT, O 
                           => G_4350GAT_OUT);
   G_4349GAT : Nor_gate port map( I1 => G_4290GAT_OUT, I2 => G_1248GAT_OUT, O 
                           => G_4349GAT_OUT);
   G_4348GAT : Nor_gate port map( I1 => G_4238GAT_OUT, I2 => G_4290GAT_OUT, O 
                           => G_4348GAT_OUT);
   G_4344GAT : Nor_gate port map( I1 => G_4287GAT_OUT, I2 => G_1200GAT_OUT, O 
                           => G_4344GAT_OUT);
   G_4341GAT : Nor_gate port map( I1 => G_4285GAT_OUT, I2 => G_4286GAT_OUT, O 
                           => G_4341GAT_OUT);
   G_4340GAT : Nor_gate port map( I1 => G_4281GAT_OUT, I2 => G_4226GAT_OUT, O 
                           => G_4340GAT_OUT);
   G_4339GAT : Nor_gate port map( I1 => G_4229GAT_OUT, I2 => G_4281GAT_OUT, O 
                           => G_4339GAT_OUT);
   G_4335GAT : Nor_gate port map( I1 => G_4278GAT_OUT, I2 => G_4275GAT_OUT, O 
                           => G_4335GAT_OUT);
   G_4332GAT : Nor_gate port map( I1 => G_4273GAT_OUT, I2 => G_4274GAT_OUT, O 
                           => G_4332GAT_OUT);
   G_4329GAT : Nor_gate port map( I1 => G_4085GAT_OUT, I2 => G_4269GAT_OUT, O 
                           => G_4329GAT_OUT);
   G_4328GAT : Nor_gate port map( I1 => G_4269GAT_OUT, I2 => G_1005GAT_OUT, O 
                           => G_4328GAT_OUT);
   G_4327GAT : Nor_gate port map( I1 => G_4217GAT_OUT, I2 => G_4269GAT_OUT, O 
                           => G_4327GAT_OUT);
   G_4323GAT : Nor_gate port map( I1 => G_4266GAT_OUT, I2 => G_957GAT_OUT, O =>
                           G_4323GAT_OUT);
   G_4320GAT : Nor_gate port map( I1 => G_4264GAT_OUT, I2 => G_4265GAT_OUT, O 
                           => G_4320GAT_OUT);
   G_4319GAT : Nor_gate port map( I1 => G_4260GAT_OUT, I2 => G_4205GAT_OUT, O 
                           => G_4319GAT_OUT);
   G_4318GAT : Nor_gate port map( I1 => G_4208GAT_OUT, I2 => G_4260GAT_OUT, O 
                           => G_4318GAT_OUT);
   G_4314GAT : Nor_gate port map( I1 => G_4257GAT_OUT, I2 => G_4200GAT_OUT, O 
                           => G_4314GAT_OUT);
   G_4310GAT : Nor_gate port map( I1 => G_4254GAT_OUT, I2 => G_4195GAT_OUT, O 
                           => G_4310GAT_OUT);
   G_4306GAT : Nor_gate port map( I1 => G_4251GAT_OUT, I2 => G_4190GAT_OUT, O 
                           => G_4306GAT_OUT);
   G_4302GAT : Nor_gate port map( I1 => G_4248GAT_OUT, I2 => G_4185GAT_OUT, O 
                           => G_4302GAT_OUT);
   G_4298GAT : Nor_gate port map( I1 => G_4245GAT_OUT, I2 => G_4180GAT_OUT, O 
                           => G_4298GAT_OUT);
   G_4294GAT : Nor_gate port map( I1 => G_4242GAT_OUT, I2 => G_4175GAT_OUT, O 
                           => G_4294GAT_OUT);
   G_4290GAT : Nor_gate port map( I1 => G_4238GAT_OUT, I2 => G_1248GAT_OUT, O 
                           => G_4290GAT_OUT);
   G_4287GAT : Nor_gate port map( I1 => G_4236GAT_OUT, I2 => G_4237GAT_OUT, O 
                           => G_4287GAT_OUT);
   G_4286GAT : Nor_gate port map( I1 => G_4232GAT_OUT, I2 => G_4161GAT_OUT, O 
                           => G_4286GAT_OUT);
   G_4285GAT : Nor_gate port map( I1 => G_4164GAT_OUT, I2 => G_4232GAT_OUT, O 
                           => G_4285GAT_OUT);
   G_4281GAT : Nor_gate port map( I1 => G_4229GAT_OUT, I2 => G_4226GAT_OUT, O 
                           => G_4281GAT_OUT);
   G_4278GAT : Nor_gate port map( I1 => G_4224GAT_OUT, I2 => G_4225GAT_OUT, O 
                           => G_4278GAT_OUT);
   G_4275GAT : Nor_gate port map( I1 => G_4034GAT_OUT, I2 => G_4220GAT_OUT, O 
                           => G_4275GAT_OUT);
   G_4274GAT : Nor_gate port map( I1 => G_4220GAT_OUT, I2 => G_1053GAT_OUT, O 
                           => G_4274GAT_OUT);
   G_4273GAT : Nor_gate port map( I1 => G_4152GAT_OUT, I2 => G_4220GAT_OUT, O 
                           => G_4273GAT_OUT);
   G_4269GAT : Nor_gate port map( I1 => G_4217GAT_OUT, I2 => G_1005GAT_OUT, O 
                           => G_4269GAT_OUT);
   G_4266GAT : Nor_gate port map( I1 => G_4215GAT_OUT, I2 => G_4216GAT_OUT, O 
                           => G_4266GAT_OUT);
   G_4265GAT : Nor_gate port map( I1 => G_4211GAT_OUT, I2 => G_4140GAT_OUT, O 
                           => G_4265GAT_OUT);
   G_4264GAT : Nor_gate port map( I1 => G_4143GAT_OUT, I2 => G_4211GAT_OUT, O 
                           => G_4264GAT_OUT);
   G_4260GAT : Nor_gate port map( I1 => G_4208GAT_OUT, I2 => G_4205GAT_OUT, O 
                           => G_4260GAT_OUT);
   G_4257GAT : Nor_gate port map( I1 => G_4203GAT_OUT, I2 => G_4204GAT_OUT, O 
                           => G_4257GAT_OUT);
   G_4254GAT : Nor_gate port map( I1 => G_4198GAT_OUT, I2 => G_4199GAT_OUT, O 
                           => G_4254GAT_OUT);
   G_4251GAT : Nor_gate port map( I1 => G_4193GAT_OUT, I2 => G_4194GAT_OUT, O 
                           => G_4251GAT_OUT);
   G_4248GAT : Nor_gate port map( I1 => G_4188GAT_OUT, I2 => G_4189GAT_OUT, O 
                           => G_4248GAT_OUT);
   G_4245GAT : Nor_gate port map( I1 => G_4183GAT_OUT, I2 => G_4184GAT_OUT, O 
                           => G_4245GAT_OUT);
   G_4242GAT : Nor_gate port map( I1 => G_4178GAT_OUT, I2 => G_4179GAT_OUT, O 
                           => G_4242GAT_OUT);
   G_4238GAT : Nor_gate port map( I1 => G_4171GAT_OUT, I2 => G_4172GAT_OUT, O 
                           => G_4238GAT_OUT);
   G_4237GAT : Nor_gate port map( I1 => G_4167GAT_OUT, I2 => G_4100GAT_OUT, O 
                           => G_4237GAT_OUT);
   G_4236GAT : Nor_gate port map( I1 => G_4103GAT_OUT, I2 => G_4167GAT_OUT, O 
                           => G_4236GAT_OUT);
   G_4232GAT : Nor_gate port map( I1 => G_4164GAT_OUT, I2 => G_4161GAT_OUT, O 
                           => G_4232GAT_OUT);
   G_4229GAT : Nor_gate port map( I1 => G_4159GAT_OUT, I2 => G_4160GAT_OUT, O 
                           => G_4229GAT_OUT);
   G_4226GAT : Nor_gate port map( I1 => G_3992GAT_OUT, I2 => G_4155GAT_OUT, O 
                           => G_4226GAT_OUT);
   G_4225GAT : Nor_gate port map( I1 => G_4155GAT_OUT, I2 => G_1101GAT_OUT, O 
                           => G_4225GAT_OUT);
   G_4224GAT : Nor_gate port map( I1 => G_4091GAT_OUT, I2 => G_4155GAT_OUT, O 
                           => G_4224GAT_OUT);
   G_4220GAT : Nor_gate port map( I1 => G_4152GAT_OUT, I2 => G_1053GAT_OUT, O 
                           => G_4220GAT_OUT);
   G_4217GAT : Nor_gate port map( I1 => G_4150GAT_OUT, I2 => G_4151GAT_OUT, O 
                           => G_4217GAT_OUT);
   G_4216GAT : Nor_gate port map( I1 => G_4146GAT_OUT, I2 => G_4079GAT_OUT, O 
                           => G_4216GAT_OUT);
   G_4215GAT : Nor_gate port map( I1 => G_4082GAT_OUT, I2 => G_4146GAT_OUT, O 
                           => G_4215GAT_OUT);
   G_4211GAT : Nor_gate port map( I1 => G_4143GAT_OUT, I2 => G_4140GAT_OUT, O 
                           => G_4211GAT_OUT);
   G_4208GAT : Nor_gate port map( I1 => G_4138GAT_OUT, I2 => G_4139GAT_OUT, O 
                           => G_4208GAT_OUT);
   G_4205GAT : Nor_gate port map( I1 => G_3971GAT_OUT, I2 => G_4134GAT_OUT, O 
                           => G_4205GAT_OUT);
   G_4204GAT : Nor_gate port map( I1 => G_4134GAT_OUT, I2 => G_858GAT_OUT, O =>
                           G_4204GAT_OUT);
   G_4203GAT : Nor_gate port map( I1 => G_4070GAT_OUT, I2 => G_4134GAT_OUT, O 
                           => G_4203GAT_OUT);
   G_4200GAT : Nor_gate port map( I1 => G_3967GAT_OUT, I2 => G_4130GAT_OUT, O 
                           => G_4200GAT_OUT);
   G_4199GAT : Nor_gate port map( I1 => G_4130GAT_OUT, I2 => G_810GAT_OUT, O =>
                           G_4199GAT_OUT);
   G_4198GAT : Nor_gate port map( I1 => G_4067GAT_OUT, I2 => G_4130GAT_OUT, O 
                           => G_4198GAT_OUT);
   G_4195GAT : Nor_gate port map( I1 => G_3963GAT_OUT, I2 => G_4126GAT_OUT, O 
                           => G_4195GAT_OUT);
   G_4194GAT : Nor_gate port map( I1 => G_4126GAT_OUT, I2 => G_762GAT_OUT, O =>
                           G_4194GAT_OUT);
   G_4193GAT : Nor_gate port map( I1 => G_4064GAT_OUT, I2 => G_4126GAT_OUT, O 
                           => G_4193GAT_OUT);
   G_4190GAT : Nor_gate port map( I1 => G_3959GAT_OUT, I2 => G_4122GAT_OUT, O 
                           => G_4190GAT_OUT);
   G_4189GAT : Nor_gate port map( I1 => G_4122GAT_OUT, I2 => G_714GAT_OUT, O =>
                           G_4189GAT_OUT);
   G_4188GAT : Nor_gate port map( I1 => G_4061GAT_OUT, I2 => G_4122GAT_OUT, O 
                           => G_4188GAT_OUT);
   G_4185GAT : Nor_gate port map( I1 => G_3955GAT_OUT, I2 => G_4118GAT_OUT, O 
                           => G_4185GAT_OUT);
   G_4184GAT : Nor_gate port map( I1 => G_4118GAT_OUT, I2 => G_666GAT_OUT, O =>
                           G_4184GAT_OUT);
   G_4183GAT : Nor_gate port map( I1 => G_4058GAT_OUT, I2 => G_4118GAT_OUT, O 
                           => G_4183GAT_OUT);
   G_4180GAT : Nor_gate port map( I1 => G_3951GAT_OUT, I2 => G_4114GAT_OUT, O 
                           => G_4180GAT_OUT);
   G_4179GAT : Nor_gate port map( I1 => G_4114GAT_OUT, I2 => G_618GAT_OUT, O =>
                           G_4179GAT_OUT);
   G_4178GAT : Nor_gate port map( I1 => G_4055GAT_OUT, I2 => G_4114GAT_OUT, O 
                           => G_4178GAT_OUT);
   G_4175GAT : Nor_gate port map( I1 => G_3947GAT_OUT, I2 => G_4110GAT_OUT, O 
                           => G_4175GAT_OUT);
   G_4174GAT : Nor_gate port map( I1 => G_4110GAT_OUT, I2 => G_570GAT_OUT, O =>
                           G_4174GAT_OUT);
   G_4173GAT : Nor_gate port map( I1 => G_4052GAT_OUT, I2 => G_4110GAT_OUT, O 
                           => G_4173GAT_OUT);
   G_4172GAT : Nor_gate port map( I1 => G_4106GAT_OUT, I2 => G_4049GAT_OUT, O 
                           => G_4172GAT_OUT);
   G_4171GAT : Nor_gate port map( I1 => G_1293GAT_OUT, I2 => G_4106GAT_OUT, O 
                           => G_4171GAT_OUT);
   G_4167GAT : Nor_gate port map( I1 => G_4103GAT_OUT, I2 => G_4100GAT_OUT, O 
                           => G_4167GAT_OUT);
   G_4164GAT : Nor_gate port map( I1 => G_4098GAT_OUT, I2 => G_4099GAT_OUT, O 
                           => G_4164GAT_OUT);
   G_4161GAT : Nor_gate port map( I1 => G_3938GAT_OUT, I2 => G_4094GAT_OUT, O 
                           => G_4161GAT_OUT);
   G_4160GAT : Nor_gate port map( I1 => G_4094GAT_OUT, I2 => G_1149GAT_OUT, O 
                           => G_4160GAT_OUT);
   G_4159GAT : Nor_gate port map( I1 => G_4040GAT_OUT, I2 => G_4094GAT_OUT, O 
                           => G_4159GAT_OUT);
   G_4155GAT : Nor_gate port map( I1 => G_4091GAT_OUT, I2 => G_1101GAT_OUT, O 
                           => G_4155GAT_OUT);
   G_4152GAT : Nor_gate port map( I1 => G_4089GAT_OUT, I2 => G_4090GAT_OUT, O 
                           => G_4152GAT_OUT);
   G_4151GAT : Nor_gate port map( I1 => G_4085GAT_OUT, I2 => G_4028GAT_OUT, O 
                           => G_4151GAT_OUT);
   G_4150GAT : Nor_gate port map( I1 => G_4031GAT_OUT, I2 => G_4085GAT_OUT, O 
                           => G_4150GAT_OUT);
   G_4146GAT : Nor_gate port map( I1 => G_4082GAT_OUT, I2 => G_4079GAT_OUT, O 
                           => G_4146GAT_OUT);
   G_4143GAT : Nor_gate port map( I1 => G_4077GAT_OUT, I2 => G_4078GAT_OUT, O 
                           => G_4143GAT_OUT);
   G_4140GAT : Nor_gate port map( I1 => G_3917GAT_OUT, I2 => G_4073GAT_OUT, O 
                           => G_4140GAT_OUT);
   G_4139GAT : Nor_gate port map( I1 => G_4073GAT_OUT, I2 => G_906GAT_OUT, O =>
                           G_4139GAT_OUT);
   G_4138GAT : Nor_gate port map( I1 => G_4019GAT_OUT, I2 => G_4073GAT_OUT, O 
                           => G_4138GAT_OUT);
   G_4134GAT : Nor_gate port map( I1 => G_4070GAT_OUT, I2 => G_858GAT_OUT, O =>
                           G_4134GAT_OUT);
   G_4130GAT : Nor_gate port map( I1 => G_4067GAT_OUT, I2 => G_810GAT_OUT, O =>
                           G_4130GAT_OUT);
   G_4126GAT : Nor_gate port map( I1 => G_4064GAT_OUT, I2 => G_762GAT_OUT, O =>
                           G_4126GAT_OUT);
   G_4122GAT : Nor_gate port map( I1 => G_4061GAT_OUT, I2 => G_714GAT_OUT, O =>
                           G_4122GAT_OUT);
   G_4118GAT : Nor_gate port map( I1 => G_4058GAT_OUT, I2 => G_666GAT_OUT, O =>
                           G_4118GAT_OUT);
   G_4114GAT : Nor_gate port map( I1 => G_4055GAT_OUT, I2 => G_618GAT_OUT, O =>
                           G_4114GAT_OUT);
   G_4110GAT : Nor_gate port map( I1 => G_4052GAT_OUT, I2 => G_570GAT_OUT, O =>
                           G_4110GAT_OUT);
   G_4106GAT : Nor_gate port map( I1 => G_1293GAT_OUT, I2 => G_4049GAT_OUT, O 
                           => G_4106GAT_OUT);
   G_4103GAT : Nor_gate port map( I1 => G_4047GAT_OUT, I2 => G_4048GAT_OUT, O 
                           => G_4103GAT_OUT);
   G_4100GAT : Nor_gate port map( I1 => G_3889GAT_OUT, I2 => G_4043GAT_OUT, O 
                           => G_4100GAT_OUT);
   G_4099GAT : Nor_gate port map( I1 => G_4043GAT_OUT, I2 => G_1197GAT_OUT, O 
                           => G_4099GAT_OUT);
   G_4098GAT : Nor_gate port map( I1 => G_3998GAT_OUT, I2 => G_4043GAT_OUT, O 
                           => G_4098GAT_OUT);
   G_4094GAT : Nor_gate port map( I1 => G_4040GAT_OUT, I2 => G_1149GAT_OUT, O 
                           => G_4094GAT_OUT);
   G_4091GAT : Nor_gate port map( I1 => G_4038GAT_OUT, I2 => G_4039GAT_OUT, O 
                           => G_4091GAT_OUT);
   G_4090GAT : Nor_gate port map( I1 => G_4034GAT_OUT, I2 => G_3986GAT_OUT, O 
                           => G_4090GAT_OUT);
   G_4089GAT : Nor_gate port map( I1 => G_3989GAT_OUT, I2 => G_4034GAT_OUT, O 
                           => G_4089GAT_OUT);
   G_4085GAT : Nor_gate port map( I1 => G_4031GAT_OUT, I2 => G_4028GAT_OUT, O 
                           => G_4085GAT_OUT);
   G_4082GAT : Nor_gate port map( I1 => G_4026GAT_OUT, I2 => G_4027GAT_OUT, O 
                           => G_4082GAT_OUT);
   G_4079GAT : Nor_gate port map( I1 => G_3868GAT_OUT, I2 => G_4022GAT_OUT, O 
                           => G_4079GAT_OUT);
   G_4078GAT : Nor_gate port map( I1 => G_4022GAT_OUT, I2 => G_954GAT_OUT, O =>
                           G_4078GAT_OUT);
   G_4077GAT : Nor_gate port map( I1 => G_3977GAT_OUT, I2 => G_4022GAT_OUT, O 
                           => G_4077GAT_OUT);
   G_4073GAT : Nor_gate port map( I1 => G_4019GAT_OUT, I2 => G_906GAT_OUT, O =>
                           G_4073GAT_OUT);
   G_4070GAT : Nor_gate port map( I1 => G_4017GAT_OUT, I2 => G_4018GAT_OUT, O 
                           => G_4070GAT_OUT);
   G_4067GAT : Nor_gate port map( I1 => G_4015GAT_OUT, I2 => G_4016GAT_OUT, O 
                           => G_4067GAT_OUT);
   G_4064GAT : Nor_gate port map( I1 => G_4013GAT_OUT, I2 => G_4014GAT_OUT, O 
                           => G_4064GAT_OUT);
   G_4061GAT : Nor_gate port map( I1 => G_4011GAT_OUT, I2 => G_4012GAT_OUT, O 
                           => G_4061GAT_OUT);
   G_4058GAT : Nor_gate port map( I1 => G_4009GAT_OUT, I2 => G_4010GAT_OUT, O 
                           => G_4058GAT_OUT);
   G_4055GAT : Nor_gate port map( I1 => G_4007GAT_OUT, I2 => G_4008GAT_OUT, O 
                           => G_4055GAT_OUT);
   G_4052GAT : Nor_gate port map( I1 => G_4005GAT_OUT, I2 => G_4006GAT_OUT, O 
                           => G_4052GAT_OUT);
   G_4049GAT : Nor_gate port map( I1 => G_3821GAT_OUT, I2 => G_4001GAT_OUT, O 
                           => G_4049GAT_OUT);
   G_4048GAT : Nor_gate port map( I1 => G_4001GAT_OUT, I2 => G_1245GAT_OUT, O 
                           => G_4048GAT_OUT);
   G_4047GAT : Nor_gate port map( I1 => G_3944GAT_OUT, I2 => G_4001GAT_OUT, O 
                           => G_4047GAT_OUT);
   G_4043GAT : Nor_gate port map( I1 => G_3998GAT_OUT, I2 => G_1197GAT_OUT, O 
                           => G_4043GAT_OUT);
   G_4040GAT : Nor_gate port map( I1 => G_3996GAT_OUT, I2 => G_3997GAT_OUT, O 
                           => G_4040GAT_OUT);
   G_4039GAT : Nor_gate port map( I1 => G_3992GAT_OUT, I2 => G_3932GAT_OUT, O 
                           => G_4039GAT_OUT);
   G_4038GAT : Nor_gate port map( I1 => G_3935GAT_OUT, I2 => G_3992GAT_OUT, O 
                           => G_4038GAT_OUT);
   G_4034GAT : Nor_gate port map( I1 => G_3989GAT_OUT, I2 => G_3986GAT_OUT, O 
                           => G_4034GAT_OUT);
   G_4031GAT : Nor_gate port map( I1 => G_3984GAT_OUT, I2 => G_3985GAT_OUT, O 
                           => G_4031GAT_OUT);
   G_4028GAT : Nor_gate port map( I1 => G_3800GAT_OUT, I2 => G_3980GAT_OUT, O 
                           => G_4028GAT_OUT);
   G_4027GAT : Nor_gate port map( I1 => G_3980GAT_OUT, I2 => G_1002GAT_OUT, O 
                           => G_4027GAT_OUT);
   G_4026GAT : Nor_gate port map( I1 => G_3923GAT_OUT, I2 => G_3980GAT_OUT, O 
                           => G_4026GAT_OUT);
   G_4022GAT : Nor_gate port map( I1 => G_3977GAT_OUT, I2 => G_954GAT_OUT, O =>
                           G_4022GAT_OUT);
   G_4019GAT : Nor_gate port map( I1 => G_3975GAT_OUT, I2 => G_3976GAT_OUT, O 
                           => G_4019GAT_OUT);
   G_4018GAT : Nor_gate port map( I1 => G_3971GAT_OUT, I2 => G_3857GAT_OUT, O 
                           => G_4018GAT_OUT);
   G_4017GAT : Nor_gate port map( I1 => G_3914GAT_OUT, I2 => G_3971GAT_OUT, O 
                           => G_4017GAT_OUT);
   G_4016GAT : Nor_gate port map( I1 => G_3967GAT_OUT, I2 => G_3852GAT_OUT, O 
                           => G_4016GAT_OUT);
   G_4015GAT : Nor_gate port map( I1 => G_3911GAT_OUT, I2 => G_3967GAT_OUT, O 
                           => G_4015GAT_OUT);
   G_4014GAT : Nor_gate port map( I1 => G_3963GAT_OUT, I2 => G_3847GAT_OUT, O 
                           => G_4014GAT_OUT);
   G_4013GAT : Nor_gate port map( I1 => G_3908GAT_OUT, I2 => G_3963GAT_OUT, O 
                           => G_4013GAT_OUT);
   G_4012GAT : Nor_gate port map( I1 => G_3959GAT_OUT, I2 => G_3842GAT_OUT, O 
                           => G_4012GAT_OUT);
   G_4011GAT : Nor_gate port map( I1 => G_3905GAT_OUT, I2 => G_3959GAT_OUT, O 
                           => G_4011GAT_OUT);
   G_4010GAT : Nor_gate port map( I1 => G_3955GAT_OUT, I2 => G_3837GAT_OUT, O 
                           => G_4010GAT_OUT);
   G_4009GAT : Nor_gate port map( I1 => G_3902GAT_OUT, I2 => G_3955GAT_OUT, O 
                           => G_4009GAT_OUT);
   G_4008GAT : Nor_gate port map( I1 => G_3951GAT_OUT, I2 => G_3832GAT_OUT, O 
                           => G_4008GAT_OUT);
   G_4007GAT : Nor_gate port map( I1 => G_3899GAT_OUT, I2 => G_3951GAT_OUT, O 
                           => G_4007GAT_OUT);
   G_4006GAT : Nor_gate port map( I1 => G_3947GAT_OUT, I2 => G_3827GAT_OUT, O 
                           => G_4006GAT_OUT);
   G_4005GAT : Nor_gate port map( I1 => G_3896GAT_OUT, I2 => G_3947GAT_OUT, O 
                           => G_4005GAT_OUT);
   G_4001GAT : Nor_gate port map( I1 => G_3944GAT_OUT, I2 => G_1245GAT_OUT, O 
                           => G_4001GAT_OUT);
   G_3998GAT : Nor_gate port map( I1 => G_3942GAT_OUT, I2 => G_3943GAT_OUT, O 
                           => G_3998GAT_OUT);
   G_3997GAT : Nor_gate port map( I1 => G_3938GAT_OUT, I2 => G_3883GAT_OUT, O 
                           => G_3997GAT_OUT);
   G_3996GAT : Nor_gate port map( I1 => G_3886GAT_OUT, I2 => G_3938GAT_OUT, O 
                           => G_3996GAT_OUT);
   G_3992GAT : Nor_gate port map( I1 => G_3935GAT_OUT, I2 => G_3932GAT_OUT, O 
                           => G_3992GAT_OUT);
   G_3989GAT : Nor_gate port map( I1 => G_3930GAT_OUT, I2 => G_3931GAT_OUT, O 
                           => G_3989GAT_OUT);
   G_3986GAT : Nor_gate port map( I1 => G_3742GAT_OUT, I2 => G_3926GAT_OUT, O 
                           => G_3986GAT_OUT);
   G_3985GAT : Nor_gate port map( I1 => G_3926GAT_OUT, I2 => G_1050GAT_OUT, O 
                           => G_3985GAT_OUT);
   G_3984GAT : Nor_gate port map( I1 => G_3874GAT_OUT, I2 => G_3926GAT_OUT, O 
                           => G_3984GAT_OUT);
   G_3980GAT : Nor_gate port map( I1 => G_3923GAT_OUT, I2 => G_1002GAT_OUT, O 
                           => G_3980GAT_OUT);
   G_3977GAT : Nor_gate port map( I1 => G_3921GAT_OUT, I2 => G_3922GAT_OUT, O 
                           => G_3977GAT_OUT);
   G_3976GAT : Nor_gate port map( I1 => G_3917GAT_OUT, I2 => G_3862GAT_OUT, O 
                           => G_3976GAT_OUT);
   G_3975GAT : Nor_gate port map( I1 => G_3865GAT_OUT, I2 => G_3917GAT_OUT, O 
                           => G_3975GAT_OUT);
   G_3971GAT : Nor_gate port map( I1 => G_3914GAT_OUT, I2 => G_3857GAT_OUT, O 
                           => G_3971GAT_OUT);
   G_3967GAT : Nor_gate port map( I1 => G_3911GAT_OUT, I2 => G_3852GAT_OUT, O 
                           => G_3967GAT_OUT);
   G_3963GAT : Nor_gate port map( I1 => G_3908GAT_OUT, I2 => G_3847GAT_OUT, O 
                           => G_3963GAT_OUT);
   G_3959GAT : Nor_gate port map( I1 => G_3905GAT_OUT, I2 => G_3842GAT_OUT, O 
                           => G_3959GAT_OUT);
   G_3955GAT : Nor_gate port map( I1 => G_3902GAT_OUT, I2 => G_3837GAT_OUT, O 
                           => G_3955GAT_OUT);
   G_3951GAT : Nor_gate port map( I1 => G_3899GAT_OUT, I2 => G_3832GAT_OUT, O 
                           => G_3951GAT_OUT);
   G_3947GAT : Nor_gate port map( I1 => G_3896GAT_OUT, I2 => G_3827GAT_OUT, O 
                           => G_3947GAT_OUT);
   G_3944GAT : Nor_gate port map( I1 => G_3893GAT_OUT, I2 => G_3894GAT_OUT, O 
                           => G_3944GAT_OUT);
   G_3943GAT : Nor_gate port map( I1 => G_3889GAT_OUT, I2 => G_3815GAT_OUT, O 
                           => G_3943GAT_OUT);
   G_3942GAT : Nor_gate port map( I1 => G_3818GAT_OUT, I2 => G_3889GAT_OUT, O 
                           => G_3942GAT_OUT);
   G_3938GAT : Nor_gate port map( I1 => G_3886GAT_OUT, I2 => G_3883GAT_OUT, O 
                           => G_3938GAT_OUT);
   G_3935GAT : Nor_gate port map( I1 => G_3881GAT_OUT, I2 => G_3882GAT_OUT, O 
                           => G_3935GAT_OUT);
   G_3932GAT : Nor_gate port map( I1 => G_3693GAT_OUT, I2 => G_3877GAT_OUT, O 
                           => G_3932GAT_OUT);
   G_3931GAT : Nor_gate port map( I1 => G_3877GAT_OUT, I2 => G_1098GAT_OUT, O 
                           => G_3931GAT_OUT);
   G_3930GAT : Nor_gate port map( I1 => G_3806GAT_OUT, I2 => G_3877GAT_OUT, O 
                           => G_3930GAT_OUT);
   G_3926GAT : Nor_gate port map( I1 => G_3874GAT_OUT, I2 => G_1050GAT_OUT, O 
                           => G_3926GAT_OUT);
   G_3923GAT : Nor_gate port map( I1 => G_3872GAT_OUT, I2 => G_3873GAT_OUT, O 
                           => G_3923GAT_OUT);
   G_3922GAT : Nor_gate port map( I1 => G_3868GAT_OUT, I2 => G_3794GAT_OUT, O 
                           => G_3922GAT_OUT);
   G_3921GAT : Nor_gate port map( I1 => G_3797GAT_OUT, I2 => G_3868GAT_OUT, O 
                           => G_3921GAT_OUT);
   G_3917GAT : Nor_gate port map( I1 => G_3865GAT_OUT, I2 => G_3862GAT_OUT, O 
                           => G_3917GAT_OUT);
   G_3914GAT : Nor_gate port map( I1 => G_3860GAT_OUT, I2 => G_3861GAT_OUT, O 
                           => G_3914GAT_OUT);
   G_3911GAT : Nor_gate port map( I1 => G_3855GAT_OUT, I2 => G_3856GAT_OUT, O 
                           => G_3911GAT_OUT);
   G_3908GAT : Nor_gate port map( I1 => G_3850GAT_OUT, I2 => G_3851GAT_OUT, O 
                           => G_3908GAT_OUT);
   G_3905GAT : Nor_gate port map( I1 => G_3845GAT_OUT, I2 => G_3846GAT_OUT, O 
                           => G_3905GAT_OUT);
   G_3902GAT : Nor_gate port map( I1 => G_3840GAT_OUT, I2 => G_3841GAT_OUT, O 
                           => G_3902GAT_OUT);
   G_3899GAT : Nor_gate port map( I1 => G_3835GAT_OUT, I2 => G_3836GAT_OUT, O 
                           => G_3899GAT_OUT);
   G_3896GAT : Nor_gate port map( I1 => G_3830GAT_OUT, I2 => G_3831GAT_OUT, O 
                           => G_3896GAT_OUT);
   G_3894GAT : Nor_gate port map( I1 => G_3821GAT_OUT, I2 => G_3757GAT_OUT, O 
                           => G_3894GAT_OUT);
   G_3893GAT : Nor_gate port map( I1 => G_1290GAT_OUT, I2 => G_3821GAT_OUT, O 
                           => G_3893GAT_OUT);
   G_3889GAT : Nor_gate port map( I1 => G_3818GAT_OUT, I2 => G_3815GAT_OUT, O 
                           => G_3889GAT_OUT);
   G_3886GAT : Nor_gate port map( I1 => G_3813GAT_OUT, I2 => G_3814GAT_OUT, O 
                           => G_3886GAT_OUT);
   G_3883GAT : Nor_gate port map( I1 => G_3653GAT_OUT, I2 => G_3809GAT_OUT, O 
                           => G_3883GAT_OUT);
   G_3882GAT : Nor_gate port map( I1 => G_3809GAT_OUT, I2 => G_1146GAT_OUT, O 
                           => G_3882GAT_OUT);
   G_3881GAT : Nor_gate port map( I1 => G_3748GAT_OUT, I2 => G_3809GAT_OUT, O 
                           => G_3881GAT_OUT);
   G_3877GAT : Nor_gate port map( I1 => G_3806GAT_OUT, I2 => G_1098GAT_OUT, O 
                           => G_3877GAT_OUT);
   G_3874GAT : Nor_gate port map( I1 => G_3804GAT_OUT, I2 => G_3805GAT_OUT, O 
                           => G_3874GAT_OUT);
   G_3873GAT : Nor_gate port map( I1 => G_3800GAT_OUT, I2 => G_3736GAT_OUT, O 
                           => G_3873GAT_OUT);
   G_3872GAT : Nor_gate port map( I1 => G_3739GAT_OUT, I2 => G_3800GAT_OUT, O 
                           => G_3872GAT_OUT);
   G_3868GAT : Nor_gate port map( I1 => G_3797GAT_OUT, I2 => G_3794GAT_OUT, O 
                           => G_3868GAT_OUT);
   G_3865GAT : Nor_gate port map( I1 => G_3792GAT_OUT, I2 => G_3793GAT_OUT, O 
                           => G_3865GAT_OUT);
   G_3862GAT : Nor_gate port map( I1 => G_3632GAT_OUT, I2 => G_3788GAT_OUT, O 
                           => G_3862GAT_OUT);
   G_3861GAT : Nor_gate port map( I1 => G_3788GAT_OUT, I2 => G_903GAT_OUT, O =>
                           G_3861GAT_OUT);
   G_3860GAT : Nor_gate port map( I1 => G_3727GAT_OUT, I2 => G_3788GAT_OUT, O 
                           => G_3860GAT_OUT);
   G_3857GAT : Nor_gate port map( I1 => G_3628GAT_OUT, I2 => G_3784GAT_OUT, O 
                           => G_3857GAT_OUT);
   G_3856GAT : Nor_gate port map( I1 => G_3784GAT_OUT, I2 => G_855GAT_OUT, O =>
                           G_3856GAT_OUT);
   G_3855GAT : Nor_gate port map( I1 => G_3724GAT_OUT, I2 => G_3784GAT_OUT, O 
                           => G_3855GAT_OUT);
   G_3852GAT : Nor_gate port map( I1 => G_3624GAT_OUT, I2 => G_3780GAT_OUT, O 
                           => G_3852GAT_OUT);
   G_3851GAT : Nor_gate port map( I1 => G_3780GAT_OUT, I2 => G_807GAT_OUT, O =>
                           G_3851GAT_OUT);
   G_3850GAT : Nor_gate port map( I1 => G_3721GAT_OUT, I2 => G_3780GAT_OUT, O 
                           => G_3850GAT_OUT);
   G_3847GAT : Nor_gate port map( I1 => G_3620GAT_OUT, I2 => G_3776GAT_OUT, O 
                           => G_3847GAT_OUT);
   G_3846GAT : Nor_gate port map( I1 => G_3776GAT_OUT, I2 => G_759GAT_OUT, O =>
                           G_3846GAT_OUT);
   G_3845GAT : Nor_gate port map( I1 => G_3718GAT_OUT, I2 => G_3776GAT_OUT, O 
                           => G_3845GAT_OUT);
   G_3842GAT : Nor_gate port map( I1 => G_3616GAT_OUT, I2 => G_3772GAT_OUT, O 
                           => G_3842GAT_OUT);
   G_3841GAT : Nor_gate port map( I1 => G_3772GAT_OUT, I2 => G_711GAT_OUT, O =>
                           G_3841GAT_OUT);
   G_3840GAT : Nor_gate port map( I1 => G_3715GAT_OUT, I2 => G_3772GAT_OUT, O 
                           => G_3840GAT_OUT);
   G_3837GAT : Nor_gate port map( I1 => G_3612GAT_OUT, I2 => G_3768GAT_OUT, O 
                           => G_3837GAT_OUT);
   G_3836GAT : Nor_gate port map( I1 => G_3768GAT_OUT, I2 => G_663GAT_OUT, O =>
                           G_3836GAT_OUT);
   G_3835GAT : Nor_gate port map( I1 => G_3712GAT_OUT, I2 => G_3768GAT_OUT, O 
                           => G_3835GAT_OUT);
   G_3832GAT : Nor_gate port map( I1 => G_3608GAT_OUT, I2 => G_3764GAT_OUT, O 
                           => G_3832GAT_OUT);
   G_3831GAT : Nor_gate port map( I1 => G_3764GAT_OUT, I2 => G_615GAT_OUT, O =>
                           G_3831GAT_OUT);
   G_3830GAT : Nor_gate port map( I1 => G_3709GAT_OUT, I2 => G_3764GAT_OUT, O 
                           => G_3830GAT_OUT);
   G_3827GAT : Nor_gate port map( I1 => G_3604GAT_OUT, I2 => G_3760GAT_OUT, O 
                           => G_3827GAT_OUT);
   G_3826GAT : Nor_gate port map( I1 => G_3760GAT_OUT, I2 => G_567GAT_OUT, O =>
                           G_3826GAT_OUT);
   G_3825GAT : Nor_gate port map( I1 => G_3706GAT_OUT, I2 => G_3760GAT_OUT, O 
                           => G_3825GAT_OUT);
   G_3821GAT : Nor_gate port map( I1 => G_1290GAT_OUT, I2 => G_3757GAT_OUT, O 
                           => G_3821GAT_OUT);
   G_3818GAT : Nor_gate port map( I1 => G_3755GAT_OUT, I2 => G_3756GAT_OUT, O 
                           => G_3818GAT_OUT);
   G_3815GAT : Nor_gate port map( I1 => G_3598GAT_OUT, I2 => G_3751GAT_OUT, O 
                           => G_3815GAT_OUT);
   G_3814GAT : Nor_gate port map( I1 => G_3751GAT_OUT, I2 => G_1194GAT_OUT, O 
                           => G_3814GAT_OUT);
   G_3813GAT : Nor_gate port map( I1 => G_3699GAT_OUT, I2 => G_3751GAT_OUT, O 
                           => G_3813GAT_OUT);
   G_3809GAT : Nor_gate port map( I1 => G_3748GAT_OUT, I2 => G_1146GAT_OUT, O 
                           => G_3809GAT_OUT);
   G_3806GAT : Nor_gate port map( I1 => G_3746GAT_OUT, I2 => G_3747GAT_OUT, O 
                           => G_3806GAT_OUT);
   G_3805GAT : Nor_gate port map( I1 => G_3742GAT_OUT, I2 => G_3687GAT_OUT, O 
                           => G_3805GAT_OUT);
   G_3804GAT : Nor_gate port map( I1 => G_3690GAT_OUT, I2 => G_3742GAT_OUT, O 
                           => G_3804GAT_OUT);
   G_3800GAT : Nor_gate port map( I1 => G_3739GAT_OUT, I2 => G_3736GAT_OUT, O 
                           => G_3800GAT_OUT);
   G_3797GAT : Nor_gate port map( I1 => G_3734GAT_OUT, I2 => G_3735GAT_OUT, O 
                           => G_3797GAT_OUT);
   G_3794GAT : Nor_gate port map( I1 => G_3577GAT_OUT, I2 => G_3730GAT_OUT, O 
                           => G_3794GAT_OUT);
   G_3793GAT : Nor_gate port map( I1 => G_3730GAT_OUT, I2 => G_951GAT_OUT, O =>
                           G_3793GAT_OUT);
   G_3792GAT : Nor_gate port map( I1 => G_3678GAT_OUT, I2 => G_3730GAT_OUT, O 
                           => G_3792GAT_OUT);
   G_3788GAT : Nor_gate port map( I1 => G_3727GAT_OUT, I2 => G_903GAT_OUT, O =>
                           G_3788GAT_OUT);
   G_3784GAT : Nor_gate port map( I1 => G_3724GAT_OUT, I2 => G_855GAT_OUT, O =>
                           G_3784GAT_OUT);
   G_3780GAT : Nor_gate port map( I1 => G_3721GAT_OUT, I2 => G_807GAT_OUT, O =>
                           G_3780GAT_OUT);
   G_3776GAT : Nor_gate port map( I1 => G_3718GAT_OUT, I2 => G_759GAT_OUT, O =>
                           G_3776GAT_OUT);
   G_3772GAT : Nor_gate port map( I1 => G_3715GAT_OUT, I2 => G_711GAT_OUT, O =>
                           G_3772GAT_OUT);
   G_3768GAT : Nor_gate port map( I1 => G_3712GAT_OUT, I2 => G_663GAT_OUT, O =>
                           G_3768GAT_OUT);
   G_3764GAT : Nor_gate port map( I1 => G_3709GAT_OUT, I2 => G_615GAT_OUT, O =>
                           G_3764GAT_OUT);
   G_3760GAT : Nor_gate port map( I1 => G_3706GAT_OUT, I2 => G_567GAT_OUT, O =>
                           G_3760GAT_OUT);
   G_3757GAT : Nor_gate port map( I1 => G_3548GAT_OUT, I2 => G_3702GAT_OUT, O 
                           => G_3757GAT_OUT);
   G_3756GAT : Nor_gate port map( I1 => G_3702GAT_OUT, I2 => G_1242GAT_OUT, O 
                           => G_3756GAT_OUT);
   G_3755GAT : Nor_gate port map( I1 => G_3659GAT_OUT, I2 => G_3702GAT_OUT, O 
                           => G_3755GAT_OUT);
   G_3751GAT : Nor_gate port map( I1 => G_3699GAT_OUT, I2 => G_1194GAT_OUT, O 
                           => G_3751GAT_OUT);
   G_3748GAT : Nor_gate port map( I1 => G_3697GAT_OUT, I2 => G_3698GAT_OUT, O 
                           => G_3748GAT_OUT);
   G_3747GAT : Nor_gate port map( I1 => G_3693GAT_OUT, I2 => G_3647GAT_OUT, O 
                           => G_3747GAT_OUT);
   G_3746GAT : Nor_gate port map( I1 => G_3650GAT_OUT, I2 => G_3693GAT_OUT, O 
                           => G_3746GAT_OUT);
   G_3742GAT : Nor_gate port map( I1 => G_3690GAT_OUT, I2 => G_3687GAT_OUT, O 
                           => G_3742GAT_OUT);
   G_3739GAT : Nor_gate port map( I1 => G_3685GAT_OUT, I2 => G_3686GAT_OUT, O 
                           => G_3739GAT_OUT);
   G_3736GAT : Nor_gate port map( I1 => G_3527GAT_OUT, I2 => G_3681GAT_OUT, O 
                           => G_3736GAT_OUT);
   G_3735GAT : Nor_gate port map( I1 => G_3681GAT_OUT, I2 => G_999GAT_OUT, O =>
                           G_3735GAT_OUT);
   G_3734GAT : Nor_gate port map( I1 => G_3638GAT_OUT, I2 => G_3681GAT_OUT, O 
                           => G_3734GAT_OUT);
   G_3730GAT : Nor_gate port map( I1 => G_3678GAT_OUT, I2 => G_951GAT_OUT, O =>
                           G_3730GAT_OUT);
   G_3727GAT : Nor_gate port map( I1 => G_3676GAT_OUT, I2 => G_3677GAT_OUT, O 
                           => G_3727GAT_OUT);
   G_3724GAT : Nor_gate port map( I1 => G_3674GAT_OUT, I2 => G_3675GAT_OUT, O 
                           => G_3724GAT_OUT);
   G_3721GAT : Nor_gate port map( I1 => G_3672GAT_OUT, I2 => G_3673GAT_OUT, O 
                           => G_3721GAT_OUT);
   G_3718GAT : Nor_gate port map( I1 => G_3670GAT_OUT, I2 => G_3671GAT_OUT, O 
                           => G_3718GAT_OUT);
   G_3715GAT : Nor_gate port map( I1 => G_3668GAT_OUT, I2 => G_3669GAT_OUT, O 
                           => G_3715GAT_OUT);
   G_3712GAT : Nor_gate port map( I1 => G_3666GAT_OUT, I2 => G_3667GAT_OUT, O 
                           => G_3712GAT_OUT);
   G_3709GAT : Nor_gate port map( I1 => G_3664GAT_OUT, I2 => G_3665GAT_OUT, O 
                           => G_3709GAT_OUT);
   G_3706GAT : Nor_gate port map( I1 => G_3662GAT_OUT, I2 => G_3663GAT_OUT, O 
                           => G_3706GAT_OUT);
   G_3702GAT : Nor_gate port map( I1 => G_3659GAT_OUT, I2 => G_1242GAT_OUT, O 
                           => G_3702GAT_OUT);
   G_3699GAT : Nor_gate port map( I1 => G_3657GAT_OUT, I2 => G_3658GAT_OUT, O 
                           => G_3699GAT_OUT);
   G_3698GAT : Nor_gate port map( I1 => G_3653GAT_OUT, I2 => G_3592GAT_OUT, O 
                           => G_3698GAT_OUT);
   G_3697GAT : Nor_gate port map( I1 => G_3595GAT_OUT, I2 => G_3653GAT_OUT, O 
                           => G_3697GAT_OUT);
   G_3693GAT : Nor_gate port map( I1 => G_3650GAT_OUT, I2 => G_3647GAT_OUT, O 
                           => G_3693GAT_OUT);
   G_3690GAT : Nor_gate port map( I1 => G_3645GAT_OUT, I2 => G_3646GAT_OUT, O 
                           => G_3690GAT_OUT);
   G_3687GAT : Nor_gate port map( I1 => G_3461GAT_OUT, I2 => G_3641GAT_OUT, O 
                           => G_3687GAT_OUT);
   G_3686GAT : Nor_gate port map( I1 => G_3641GAT_OUT, I2 => G_1047GAT_OUT, O 
                           => G_3686GAT_OUT);
   G_3685GAT : Nor_gate port map( I1 => G_3583GAT_OUT, I2 => G_3641GAT_OUT, O 
                           => G_3685GAT_OUT);
   G_3681GAT : Nor_gate port map( I1 => G_3638GAT_OUT, I2 => G_999GAT_OUT, O =>
                           G_3681GAT_OUT);
   G_3678GAT : Nor_gate port map( I1 => G_3636GAT_OUT, I2 => G_3637GAT_OUT, O 
                           => G_3678GAT_OUT);
   G_3677GAT : Nor_gate port map( I1 => G_3632GAT_OUT, I2 => G_3516GAT_OUT, O 
                           => G_3677GAT_OUT);
   G_3676GAT : Nor_gate port map( I1 => G_3574GAT_OUT, I2 => G_3632GAT_OUT, O 
                           => G_3676GAT_OUT);
   G_3675GAT : Nor_gate port map( I1 => G_3628GAT_OUT, I2 => G_3511GAT_OUT, O 
                           => G_3675GAT_OUT);
   G_3674GAT : Nor_gate port map( I1 => G_3571GAT_OUT, I2 => G_3628GAT_OUT, O 
                           => G_3674GAT_OUT);
   G_3673GAT : Nor_gate port map( I1 => G_3624GAT_OUT, I2 => G_3506GAT_OUT, O 
                           => G_3673GAT_OUT);
   G_3672GAT : Nor_gate port map( I1 => G_3568GAT_OUT, I2 => G_3624GAT_OUT, O 
                           => G_3672GAT_OUT);
   G_3671GAT : Nor_gate port map( I1 => G_3620GAT_OUT, I2 => G_3501GAT_OUT, O 
                           => G_3671GAT_OUT);
   G_3670GAT : Nor_gate port map( I1 => G_3565GAT_OUT, I2 => G_3620GAT_OUT, O 
                           => G_3670GAT_OUT);
   G_3669GAT : Nor_gate port map( I1 => G_3616GAT_OUT, I2 => G_3496GAT_OUT, O 
                           => G_3669GAT_OUT);
   G_3668GAT : Nor_gate port map( I1 => G_3562GAT_OUT, I2 => G_3616GAT_OUT, O 
                           => G_3668GAT_OUT);
   G_3667GAT : Nor_gate port map( I1 => G_3612GAT_OUT, I2 => G_3491GAT_OUT, O 
                           => G_3667GAT_OUT);
   G_3666GAT : Nor_gate port map( I1 => G_3559GAT_OUT, I2 => G_3612GAT_OUT, O 
                           => G_3666GAT_OUT);
   G_3665GAT : Nor_gate port map( I1 => G_3608GAT_OUT, I2 => G_3486GAT_OUT, O 
                           => G_3665GAT_OUT);
   G_3664GAT : Nor_gate port map( I1 => G_3556GAT_OUT, I2 => G_3608GAT_OUT, O 
                           => G_3664GAT_OUT);
   G_3663GAT : Nor_gate port map( I1 => G_3604GAT_OUT, I2 => G_3481GAT_OUT, O 
                           => G_3663GAT_OUT);
   G_3662GAT : Nor_gate port map( I1 => G_3553GAT_OUT, I2 => G_3604GAT_OUT, O 
                           => G_3662GAT_OUT);
   G_3659GAT : Nor_gate port map( I1 => G_3602GAT_OUT, I2 => G_3603GAT_OUT, O 
                           => G_3659GAT_OUT);
   G_3658GAT : Nor_gate port map( I1 => G_3598GAT_OUT, I2 => G_3542GAT_OUT, O 
                           => G_3658GAT_OUT);
   G_3657GAT : Nor_gate port map( I1 => G_3545GAT_OUT, I2 => G_3598GAT_OUT, O 
                           => G_3657GAT_OUT);
   G_3653GAT : Nor_gate port map( I1 => G_3595GAT_OUT, I2 => G_3592GAT_OUT, O 
                           => G_3653GAT_OUT);
   G_3650GAT : Nor_gate port map( I1 => G_3590GAT_OUT, I2 => G_3591GAT_OUT, O 
                           => G_3650GAT_OUT);
   G_3647GAT : Nor_gate port map( I1 => G_3404GAT_OUT, I2 => G_3586GAT_OUT, O 
                           => G_3647GAT_OUT);
   G_3646GAT : Nor_gate port map( I1 => G_3586GAT_OUT, I2 => G_1095GAT_OUT, O 
                           => G_3646GAT_OUT);
   G_3645GAT : Nor_gate port map( I1 => G_3533GAT_OUT, I2 => G_3586GAT_OUT, O 
                           => G_3645GAT_OUT);
   G_3641GAT : Nor_gate port map( I1 => G_3583GAT_OUT, I2 => G_1047GAT_OUT, O 
                           => G_3641GAT_OUT);
   G_3638GAT : Nor_gate port map( I1 => G_3581GAT_OUT, I2 => G_3582GAT_OUT, O 
                           => G_3638GAT_OUT);
   G_3637GAT : Nor_gate port map( I1 => G_3577GAT_OUT, I2 => G_3521GAT_OUT, O 
                           => G_3637GAT_OUT);
   G_3636GAT : Nor_gate port map( I1 => G_3524GAT_OUT, I2 => G_3577GAT_OUT, O 
                           => G_3636GAT_OUT);
   G_3632GAT : Nor_gate port map( I1 => G_3574GAT_OUT, I2 => G_3516GAT_OUT, O 
                           => G_3632GAT_OUT);
   G_3628GAT : Nor_gate port map( I1 => G_3571GAT_OUT, I2 => G_3511GAT_OUT, O 
                           => G_3628GAT_OUT);
   G_3624GAT : Nor_gate port map( I1 => G_3568GAT_OUT, I2 => G_3506GAT_OUT, O 
                           => G_3624GAT_OUT);
   G_3620GAT : Nor_gate port map( I1 => G_3565GAT_OUT, I2 => G_3501GAT_OUT, O 
                           => G_3620GAT_OUT);
   G_3616GAT : Nor_gate port map( I1 => G_3562GAT_OUT, I2 => G_3496GAT_OUT, O 
                           => G_3616GAT_OUT);
   G_3612GAT : Nor_gate port map( I1 => G_3559GAT_OUT, I2 => G_3491GAT_OUT, O 
                           => G_3612GAT_OUT);
   G_3608GAT : Nor_gate port map( I1 => G_3556GAT_OUT, I2 => G_3486GAT_OUT, O 
                           => G_3608GAT_OUT);
   G_3604GAT : Nor_gate port map( I1 => G_3553GAT_OUT, I2 => G_3481GAT_OUT, O 
                           => G_3604GAT_OUT);
   G_3603GAT : Nor_gate port map( I1 => G_3548GAT_OUT, I2 => G_3476GAT_OUT, O 
                           => G_3603GAT_OUT);
   G_3602GAT : Nor_gate port map( I1 => G_1287GAT_OUT, I2 => G_3548GAT_OUT, O 
                           => G_3602GAT_OUT);
   G_3598GAT : Nor_gate port map( I1 => G_3545GAT_OUT, I2 => G_3542GAT_OUT, O 
                           => G_3598GAT_OUT);
   G_3595GAT : Nor_gate port map( I1 => G_3540GAT_OUT, I2 => G_3541GAT_OUT, O 
                           => G_3595GAT_OUT);
   G_3592GAT : Nor_gate port map( I1 => G_3356GAT_OUT, I2 => G_3536GAT_OUT, O 
                           => G_3592GAT_OUT);
   G_3591GAT : Nor_gate port map( I1 => G_3536GAT_OUT, I2 => G_1143GAT_OUT, O 
                           => G_3591GAT_OUT);
   G_3590GAT : Nor_gate port map( I1 => G_3467GAT_OUT, I2 => G_3536GAT_OUT, O 
                           => G_3590GAT_OUT);
   G_3586GAT : Nor_gate port map( I1 => G_3533GAT_OUT, I2 => G_1095GAT_OUT, O 
                           => G_3586GAT_OUT);
   G_3583GAT : Nor_gate port map( I1 => G_3531GAT_OUT, I2 => G_3532GAT_OUT, O 
                           => G_3583GAT_OUT);
   G_3582GAT : Nor_gate port map( I1 => G_3527GAT_OUT, I2 => G_3455GAT_OUT, O 
                           => G_3582GAT_OUT);
   G_3581GAT : Nor_gate port map( I1 => G_3458GAT_OUT, I2 => G_3527GAT_OUT, O 
                           => G_3581GAT_OUT);
   G_3577GAT : Nor_gate port map( I1 => G_3524GAT_OUT, I2 => G_3521GAT_OUT, O 
                           => G_3577GAT_OUT);
   G_3574GAT : Nor_gate port map( I1 => G_3519GAT_OUT, I2 => G_3520GAT_OUT, O 
                           => G_3574GAT_OUT);
   G_3571GAT : Nor_gate port map( I1 => G_3514GAT_OUT, I2 => G_3515GAT_OUT, O 
                           => G_3571GAT_OUT);
   G_3568GAT : Nor_gate port map( I1 => G_3509GAT_OUT, I2 => G_3510GAT_OUT, O 
                           => G_3568GAT_OUT);
   G_3565GAT : Nor_gate port map( I1 => G_3504GAT_OUT, I2 => G_3505GAT_OUT, O 
                           => G_3565GAT_OUT);
   G_3562GAT : Nor_gate port map( I1 => G_3499GAT_OUT, I2 => G_3500GAT_OUT, O 
                           => G_3562GAT_OUT);
   G_3559GAT : Nor_gate port map( I1 => G_3494GAT_OUT, I2 => G_3495GAT_OUT, O 
                           => G_3559GAT_OUT);
   G_3556GAT : Nor_gate port map( I1 => G_3489GAT_OUT, I2 => G_3490GAT_OUT, O 
                           => G_3556GAT_OUT);
   G_3553GAT : Nor_gate port map( I1 => G_3484GAT_OUT, I2 => G_3485GAT_OUT, O 
                           => G_3553GAT_OUT);
   G_3548GAT : Nor_gate port map( I1 => G_1287GAT_OUT, I2 => G_3476GAT_OUT, O 
                           => G_3548GAT_OUT);
   G_3545GAT : Nor_gate port map( I1 => G_3474GAT_OUT, I2 => G_3475GAT_OUT, O 
                           => G_3545GAT_OUT);
   G_3542GAT : Nor_gate port map( I1 => G_3317GAT_OUT, I2 => G_3470GAT_OUT, O 
                           => G_3542GAT_OUT);
   G_3541GAT : Nor_gate port map( I1 => G_3470GAT_OUT, I2 => G_1191GAT_OUT, O 
                           => G_3541GAT_OUT);
   G_3540GAT : Nor_gate port map( I1 => G_3410GAT_OUT, I2 => G_3470GAT_OUT, O 
                           => G_3540GAT_OUT);
   G_3536GAT : Nor_gate port map( I1 => G_3467GAT_OUT, I2 => G_1143GAT_OUT, O 
                           => G_3536GAT_OUT);
   G_3533GAT : Nor_gate port map( I1 => G_3465GAT_OUT, I2 => G_3466GAT_OUT, O 
                           => G_3533GAT_OUT);
   G_3532GAT : Nor_gate port map( I1 => G_3461GAT_OUT, I2 => G_3398GAT_OUT, O 
                           => G_3532GAT_OUT);
   G_3531GAT : Nor_gate port map( I1 => G_3401GAT_OUT, I2 => G_3461GAT_OUT, O 
                           => G_3531GAT_OUT);
   G_3527GAT : Nor_gate port map( I1 => G_3458GAT_OUT, I2 => G_3455GAT_OUT, O 
                           => G_3527GAT_OUT);
   G_3524GAT : Nor_gate port map( I1 => G_3453GAT_OUT, I2 => G_3454GAT_OUT, O 
                           => G_3524GAT_OUT);
   G_3521GAT : Nor_gate port map( I1 => G_3296GAT_OUT, I2 => G_3449GAT_OUT, O 
                           => G_3521GAT_OUT);
   G_3520GAT : Nor_gate port map( I1 => G_3449GAT_OUT, I2 => G_948GAT_OUT, O =>
                           G_3520GAT_OUT);
   G_3519GAT : Nor_gate port map( I1 => G_3389GAT_OUT, I2 => G_3449GAT_OUT, O 
                           => G_3519GAT_OUT);
   G_3516GAT : Nor_gate port map( I1 => G_3292GAT_OUT, I2 => G_3445GAT_OUT, O 
                           => G_3516GAT_OUT);
   G_3515GAT : Nor_gate port map( I1 => G_3445GAT_OUT, I2 => G_900GAT_OUT, O =>
                           G_3515GAT_OUT);
   G_3514GAT : Nor_gate port map( I1 => G_3386GAT_OUT, I2 => G_3445GAT_OUT, O 
                           => G_3514GAT_OUT);
   G_3511GAT : Nor_gate port map( I1 => G_3288GAT_OUT, I2 => G_3441GAT_OUT, O 
                           => G_3511GAT_OUT);
   G_3510GAT : Nor_gate port map( I1 => G_3441GAT_OUT, I2 => G_852GAT_OUT, O =>
                           G_3510GAT_OUT);
   G_3509GAT : Nor_gate port map( I1 => G_3383GAT_OUT, I2 => G_3441GAT_OUT, O 
                           => G_3509GAT_OUT);
   G_3506GAT : Nor_gate port map( I1 => G_3284GAT_OUT, I2 => G_3437GAT_OUT, O 
                           => G_3506GAT_OUT);
   G_3505GAT : Nor_gate port map( I1 => G_3437GAT_OUT, I2 => G_804GAT_OUT, O =>
                           G_3505GAT_OUT);
   G_3504GAT : Nor_gate port map( I1 => G_3380GAT_OUT, I2 => G_3437GAT_OUT, O 
                           => G_3504GAT_OUT);
   G_3501GAT : Nor_gate port map( I1 => G_3280GAT_OUT, I2 => G_3433GAT_OUT, O 
                           => G_3501GAT_OUT);
   G_3500GAT : Nor_gate port map( I1 => G_3433GAT_OUT, I2 => G_756GAT_OUT, O =>
                           G_3500GAT_OUT);
   G_3499GAT : Nor_gate port map( I1 => G_3377GAT_OUT, I2 => G_3433GAT_OUT, O 
                           => G_3499GAT_OUT);
   G_3496GAT : Nor_gate port map( I1 => G_3276GAT_OUT, I2 => G_3429GAT_OUT, O 
                           => G_3496GAT_OUT);
   G_3495GAT : Nor_gate port map( I1 => G_3429GAT_OUT, I2 => G_708GAT_OUT, O =>
                           G_3495GAT_OUT);
   G_3494GAT : Nor_gate port map( I1 => G_3374GAT_OUT, I2 => G_3429GAT_OUT, O 
                           => G_3494GAT_OUT);
   G_3491GAT : Nor_gate port map( I1 => G_3272GAT_OUT, I2 => G_3425GAT_OUT, O 
                           => G_3491GAT_OUT);
   G_3490GAT : Nor_gate port map( I1 => G_3425GAT_OUT, I2 => G_660GAT_OUT, O =>
                           G_3490GAT_OUT);
   G_3489GAT : Nor_gate port map( I1 => G_3371GAT_OUT, I2 => G_3425GAT_OUT, O 
                           => G_3489GAT_OUT);
   G_3486GAT : Nor_gate port map( I1 => G_3268GAT_OUT, I2 => G_3421GAT_OUT, O 
                           => G_3486GAT_OUT);
   G_3485GAT : Nor_gate port map( I1 => G_3421GAT_OUT, I2 => G_612GAT_OUT, O =>
                           G_3485GAT_OUT);
   G_3484GAT : Nor_gate port map( I1 => G_3368GAT_OUT, I2 => G_3421GAT_OUT, O 
                           => G_3484GAT_OUT);
   G_3481GAT : Nor_gate port map( I1 => G_3264GAT_OUT, I2 => G_3417GAT_OUT, O 
                           => G_3481GAT_OUT);
   G_3480GAT : Nor_gate port map( I1 => G_3417GAT_OUT, I2 => G_564GAT_OUT, O =>
                           G_3480GAT_OUT);
   G_3479GAT : Nor_gate port map( I1 => G_3365GAT_OUT, I2 => G_3417GAT_OUT, O 
                           => G_3479GAT_OUT);
   G_3476GAT : Nor_gate port map( I1 => G_3260GAT_OUT, I2 => G_3413GAT_OUT, O 
                           => G_3476GAT_OUT);
   G_3475GAT : Nor_gate port map( I1 => G_3413GAT_OUT, I2 => G_1239GAT_OUT, O 
                           => G_3475GAT_OUT);
   G_3474GAT : Nor_gate port map( I1 => G_3362GAT_OUT, I2 => G_3413GAT_OUT, O 
                           => G_3474GAT_OUT);
   G_3470GAT : Nor_gate port map( I1 => G_3410GAT_OUT, I2 => G_1191GAT_OUT, O 
                           => G_3470GAT_OUT);
   G_3467GAT : Nor_gate port map( I1 => G_3408GAT_OUT, I2 => G_3409GAT_OUT, O 
                           => G_3467GAT_OUT);
   G_3466GAT : Nor_gate port map( I1 => G_3404GAT_OUT, I2 => G_3350GAT_OUT, O 
                           => G_3466GAT_OUT);
   G_3465GAT : Nor_gate port map( I1 => G_3353GAT_OUT, I2 => G_3404GAT_OUT, O 
                           => G_3465GAT_OUT);
   G_3461GAT : Nor_gate port map( I1 => G_3401GAT_OUT, I2 => G_3398GAT_OUT, O 
                           => G_3461GAT_OUT);
   G_3458GAT : Nor_gate port map( I1 => G_3396GAT_OUT, I2 => G_3397GAT_OUT, O 
                           => G_3458GAT_OUT);
   G_3455GAT : Nor_gate port map( I1 => G_3239GAT_OUT, I2 => G_3392GAT_OUT, O 
                           => G_3455GAT_OUT);
   G_3454GAT : Nor_gate port map( I1 => G_3392GAT_OUT, I2 => G_996GAT_OUT, O =>
                           G_3454GAT_OUT);
   G_3453GAT : Nor_gate port map( I1 => G_3341GAT_OUT, I2 => G_3392GAT_OUT, O 
                           => G_3453GAT_OUT);
   G_3449GAT : Nor_gate port map( I1 => G_3389GAT_OUT, I2 => G_948GAT_OUT, O =>
                           G_3449GAT_OUT);
   G_3445GAT : Nor_gate port map( I1 => G_3386GAT_OUT, I2 => G_900GAT_OUT, O =>
                           G_3445GAT_OUT);
   G_3441GAT : Nor_gate port map( I1 => G_3383GAT_OUT, I2 => G_852GAT_OUT, O =>
                           G_3441GAT_OUT);
   G_3437GAT : Nor_gate port map( I1 => G_3380GAT_OUT, I2 => G_804GAT_OUT, O =>
                           G_3437GAT_OUT);
   G_3433GAT : Nor_gate port map( I1 => G_3377GAT_OUT, I2 => G_756GAT_OUT, O =>
                           G_3433GAT_OUT);
   G_3429GAT : Nor_gate port map( I1 => G_3374GAT_OUT, I2 => G_708GAT_OUT, O =>
                           G_3429GAT_OUT);
   G_3425GAT : Nor_gate port map( I1 => G_3371GAT_OUT, I2 => G_660GAT_OUT, O =>
                           G_3425GAT_OUT);
   G_3421GAT : Nor_gate port map( I1 => G_3368GAT_OUT, I2 => G_612GAT_OUT, O =>
                           G_3421GAT_OUT);
   G_3417GAT : Nor_gate port map( I1 => G_3365GAT_OUT, I2 => G_564GAT_OUT, O =>
                           G_3417GAT_OUT);
   G_3413GAT : Nor_gate port map( I1 => G_3362GAT_OUT, I2 => G_1239GAT_OUT, O 
                           => G_3413GAT_OUT);
   G_3410GAT : Nor_gate port map( I1 => G_3360GAT_OUT, I2 => G_3361GAT_OUT, O 
                           => G_3410GAT_OUT);
   G_3409GAT : Nor_gate port map( I1 => G_3356GAT_OUT, I2 => G_3311GAT_OUT, O 
                           => G_3409GAT_OUT);
   G_3408GAT : Nor_gate port map( I1 => G_3314GAT_OUT, I2 => G_3356GAT_OUT, O 
                           => G_3408GAT_OUT);
   G_3404GAT : Nor_gate port map( I1 => G_3353GAT_OUT, I2 => G_3350GAT_OUT, O 
                           => G_3404GAT_OUT);
   G_3401GAT : Nor_gate port map( I1 => G_3348GAT_OUT, I2 => G_3349GAT_OUT, O 
                           => G_3401GAT_OUT);
   G_3398GAT : Nor_gate port map( I1 => G_3193GAT_OUT, I2 => G_3344GAT_OUT, O 
                           => G_3398GAT_OUT);
   G_3397GAT : Nor_gate port map( I1 => G_3344GAT_OUT, I2 => G_1044GAT_OUT, O 
                           => G_3397GAT_OUT);
   G_3396GAT : Nor_gate port map( I1 => G_3302GAT_OUT, I2 => G_3344GAT_OUT, O 
                           => G_3396GAT_OUT);
   G_3392GAT : Nor_gate port map( I1 => G_3341GAT_OUT, I2 => G_996GAT_OUT, O =>
                           G_3392GAT_OUT);
   G_3389GAT : Nor_gate port map( I1 => G_3339GAT_OUT, I2 => G_3340GAT_OUT, O 
                           => G_3389GAT_OUT);
   G_3386GAT : Nor_gate port map( I1 => G_3337GAT_OUT, I2 => G_3338GAT_OUT, O 
                           => G_3386GAT_OUT);
   G_3383GAT : Nor_gate port map( I1 => G_3335GAT_OUT, I2 => G_3336GAT_OUT, O 
                           => G_3383GAT_OUT);
   G_3380GAT : Nor_gate port map( I1 => G_3333GAT_OUT, I2 => G_3334GAT_OUT, O 
                           => G_3380GAT_OUT);
   G_3377GAT : Nor_gate port map( I1 => G_3331GAT_OUT, I2 => G_3332GAT_OUT, O 
                           => G_3377GAT_OUT);
   G_3374GAT : Nor_gate port map( I1 => G_3329GAT_OUT, I2 => G_3330GAT_OUT, O 
                           => G_3374GAT_OUT);
   G_3371GAT : Nor_gate port map( I1 => G_3327GAT_OUT, I2 => G_3328GAT_OUT, O 
                           => G_3371GAT_OUT);
   G_3368GAT : Nor_gate port map( I1 => G_3325GAT_OUT, I2 => G_3326GAT_OUT, O 
                           => G_3368GAT_OUT);
   G_3365GAT : Nor_gate port map( I1 => G_3323GAT_OUT, I2 => G_3324GAT_OUT, O 
                           => G_3365GAT_OUT);
   G_3362GAT : Nor_gate port map( I1 => G_3321GAT_OUT, I2 => G_3322GAT_OUT, O 
                           => G_3362GAT_OUT);
   G_3361GAT : Nor_gate port map( I1 => G_3317GAT_OUT, I2 => G_3254GAT_OUT, O 
                           => G_3361GAT_OUT);
   G_3360GAT : Nor_gate port map( I1 => G_3257GAT_OUT, I2 => G_3317GAT_OUT, O 
                           => G_3360GAT_OUT);
   G_3356GAT : Nor_gate port map( I1 => G_3314GAT_OUT, I2 => G_3311GAT_OUT, O 
                           => G_3356GAT_OUT);
   G_3353GAT : Nor_gate port map( I1 => G_3309GAT_OUT, I2 => G_3310GAT_OUT, O 
                           => G_3353GAT_OUT);
   G_3350GAT : Nor_gate port map( I1 => G_3127GAT_OUT, I2 => G_3305GAT_OUT, O 
                           => G_3350GAT_OUT);
   G_3349GAT : Nor_gate port map( I1 => G_3305GAT_OUT, I2 => G_1092GAT_OUT, O 
                           => G_3349GAT_OUT);
   G_3348GAT : Nor_gate port map( I1 => G_3245GAT_OUT, I2 => G_3305GAT_OUT, O 
                           => G_3348GAT_OUT);
   G_3344GAT : Nor_gate port map( I1 => G_3302GAT_OUT, I2 => G_1044GAT_OUT, O 
                           => G_3344GAT_OUT);
   G_3341GAT : Nor_gate port map( I1 => G_3300GAT_OUT, I2 => G_3301GAT_OUT, O 
                           => G_3341GAT_OUT);
   G_3340GAT : Nor_gate port map( I1 => G_3296GAT_OUT, I2 => G_3182GAT_OUT, O 
                           => G_3340GAT_OUT);
   G_3339GAT : Nor_gate port map( I1 => G_3236GAT_OUT, I2 => G_3296GAT_OUT, O 
                           => G_3339GAT_OUT);
   G_3338GAT : Nor_gate port map( I1 => G_3292GAT_OUT, I2 => G_3177GAT_OUT, O 
                           => G_3338GAT_OUT);
   G_3337GAT : Nor_gate port map( I1 => G_3233GAT_OUT, I2 => G_3292GAT_OUT, O 
                           => G_3337GAT_OUT);
   G_3336GAT : Nor_gate port map( I1 => G_3288GAT_OUT, I2 => G_3172GAT_OUT, O 
                           => G_3336GAT_OUT);
   G_3335GAT : Nor_gate port map( I1 => G_3230GAT_OUT, I2 => G_3288GAT_OUT, O 
                           => G_3335GAT_OUT);
   G_3334GAT : Nor_gate port map( I1 => G_3284GAT_OUT, I2 => G_3167GAT_OUT, O 
                           => G_3334GAT_OUT);
   G_3333GAT : Nor_gate port map( I1 => G_3227GAT_OUT, I2 => G_3284GAT_OUT, O 
                           => G_3333GAT_OUT);
   G_3332GAT : Nor_gate port map( I1 => G_3280GAT_OUT, I2 => G_3162GAT_OUT, O 
                           => G_3332GAT_OUT);
   G_3331GAT : Nor_gate port map( I1 => G_3224GAT_OUT, I2 => G_3280GAT_OUT, O 
                           => G_3331GAT_OUT);
   G_3330GAT : Nor_gate port map( I1 => G_3276GAT_OUT, I2 => G_3157GAT_OUT, O 
                           => G_3330GAT_OUT);
   G_3329GAT : Nor_gate port map( I1 => G_3221GAT_OUT, I2 => G_3276GAT_OUT, O 
                           => G_3329GAT_OUT);
   G_3328GAT : Nor_gate port map( I1 => G_3272GAT_OUT, I2 => G_3152GAT_OUT, O 
                           => G_3328GAT_OUT);
   G_3327GAT : Nor_gate port map( I1 => G_3218GAT_OUT, I2 => G_3272GAT_OUT, O 
                           => G_3327GAT_OUT);
   G_3326GAT : Nor_gate port map( I1 => G_3268GAT_OUT, I2 => G_3147GAT_OUT, O 
                           => G_3326GAT_OUT);
   G_3325GAT : Nor_gate port map( I1 => G_3215GAT_OUT, I2 => G_3268GAT_OUT, O 
                           => G_3325GAT_OUT);
   G_3324GAT : Nor_gate port map( I1 => G_3264GAT_OUT, I2 => G_3142GAT_OUT, O 
                           => G_3324GAT_OUT);
   G_3323GAT : Nor_gate port map( I1 => G_3212GAT_OUT, I2 => G_3264GAT_OUT, O 
                           => G_3323GAT_OUT);
   G_3322GAT : Nor_gate port map( I1 => G_3260GAT_OUT, I2 => G_3208GAT_OUT, O 
                           => G_3322GAT_OUT);
   G_3321GAT : Nor_gate port map( I1 => G_1284GAT_OUT, I2 => G_3260GAT_OUT, O 
                           => G_3321GAT_OUT);
   G_3317GAT : Nor_gate port map( I1 => G_3257GAT_OUT, I2 => G_3254GAT_OUT, O 
                           => G_3317GAT_OUT);
   G_3314GAT : Nor_gate port map( I1 => G_3252GAT_OUT, I2 => G_3253GAT_OUT, O 
                           => G_3314GAT_OUT);
   G_3311GAT : Nor_gate port map( I1 => G_3070GAT_OUT, I2 => G_3248GAT_OUT, O 
                           => G_3311GAT_OUT);
   G_3310GAT : Nor_gate port map( I1 => G_3248GAT_OUT, I2 => G_1140GAT_OUT, O 
                           => G_3310GAT_OUT);
   G_3309GAT : Nor_gate port map( I1 => G_3199GAT_OUT, I2 => G_3248GAT_OUT, O 
                           => G_3309GAT_OUT);
   G_3305GAT : Nor_gate port map( I1 => G_3245GAT_OUT, I2 => G_1092GAT_OUT, O 
                           => G_3305GAT_OUT);
   G_3302GAT : Nor_gate port map( I1 => G_3243GAT_OUT, I2 => G_3244GAT_OUT, O 
                           => G_3302GAT_OUT);
   G_3301GAT : Nor_gate port map( I1 => G_3239GAT_OUT, I2 => G_3187GAT_OUT, O 
                           => G_3301GAT_OUT);
   G_3300GAT : Nor_gate port map( I1 => G_3190GAT_OUT, I2 => G_3239GAT_OUT, O 
                           => G_3300GAT_OUT);
   G_3296GAT : Nor_gate port map( I1 => G_3236GAT_OUT, I2 => G_3182GAT_OUT, O 
                           => G_3296GAT_OUT);
   G_3292GAT : Nor_gate port map( I1 => G_3233GAT_OUT, I2 => G_3177GAT_OUT, O 
                           => G_3292GAT_OUT);
   G_3288GAT : Nor_gate port map( I1 => G_3230GAT_OUT, I2 => G_3172GAT_OUT, O 
                           => G_3288GAT_OUT);
   G_3284GAT : Nor_gate port map( I1 => G_3227GAT_OUT, I2 => G_3167GAT_OUT, O 
                           => G_3284GAT_OUT);
   G_3280GAT : Nor_gate port map( I1 => G_3224GAT_OUT, I2 => G_3162GAT_OUT, O 
                           => G_3280GAT_OUT);
   G_3276GAT : Nor_gate port map( I1 => G_3221GAT_OUT, I2 => G_3157GAT_OUT, O 
                           => G_3276GAT_OUT);
   G_3272GAT : Nor_gate port map( I1 => G_3218GAT_OUT, I2 => G_3152GAT_OUT, O 
                           => G_3272GAT_OUT);
   G_3268GAT : Nor_gate port map( I1 => G_3215GAT_OUT, I2 => G_3147GAT_OUT, O 
                           => G_3268GAT_OUT);
   G_3264GAT : Nor_gate port map( I1 => G_3212GAT_OUT, I2 => G_3142GAT_OUT, O 
                           => G_3264GAT_OUT);
   G_3260GAT : Nor_gate port map( I1 => G_1284GAT_OUT, I2 => G_3208GAT_OUT, O 
                           => G_3260GAT_OUT);
   G_3257GAT : Nor_gate port map( I1 => G_3206GAT_OUT, I2 => G_3207GAT_OUT, O 
                           => G_3257GAT_OUT);
   G_3254GAT : Nor_gate port map( I1 => G_3022GAT_OUT, I2 => G_3202GAT_OUT, O 
                           => G_3254GAT_OUT);
   G_3253GAT : Nor_gate port map( I1 => G_3202GAT_OUT, I2 => G_1188GAT_OUT, O 
                           => G_3253GAT_OUT);
   G_3252GAT : Nor_gate port map( I1 => G_3133GAT_OUT, I2 => G_3202GAT_OUT, O 
                           => G_3252GAT_OUT);
   G_3248GAT : Nor_gate port map( I1 => G_3199GAT_OUT, I2 => G_1140GAT_OUT, O 
                           => G_3248GAT_OUT);
   G_3245GAT : Nor_gate port map( I1 => G_3197GAT_OUT, I2 => G_3198GAT_OUT, O 
                           => G_3245GAT_OUT);
   G_3244GAT : Nor_gate port map( I1 => G_3193GAT_OUT, I2 => G_3121GAT_OUT, O 
                           => G_3244GAT_OUT);
   G_3243GAT : Nor_gate port map( I1 => G_3124GAT_OUT, I2 => G_3193GAT_OUT, O 
                           => G_3243GAT_OUT);
   G_3239GAT : Nor_gate port map( I1 => G_3190GAT_OUT, I2 => G_3187GAT_OUT, O 
                           => G_3239GAT_OUT);
   G_3236GAT : Nor_gate port map( I1 => G_3185GAT_OUT, I2 => G_3186GAT_OUT, O 
                           => G_3236GAT_OUT);
   G_3233GAT : Nor_gate port map( I1 => G_3180GAT_OUT, I2 => G_3181GAT_OUT, O 
                           => G_3233GAT_OUT);
   G_3230GAT : Nor_gate port map( I1 => G_3175GAT_OUT, I2 => G_3176GAT_OUT, O 
                           => G_3230GAT_OUT);
   G_3227GAT : Nor_gate port map( I1 => G_3170GAT_OUT, I2 => G_3171GAT_OUT, O 
                           => G_3227GAT_OUT);
   G_3224GAT : Nor_gate port map( I1 => G_3165GAT_OUT, I2 => G_3166GAT_OUT, O 
                           => G_3224GAT_OUT);
   G_3221GAT : Nor_gate port map( I1 => G_3160GAT_OUT, I2 => G_3161GAT_OUT, O 
                           => G_3221GAT_OUT);
   G_3218GAT : Nor_gate port map( I1 => G_3155GAT_OUT, I2 => G_3156GAT_OUT, O 
                           => G_3218GAT_OUT);
   G_3215GAT : Nor_gate port map( I1 => G_3150GAT_OUT, I2 => G_3151GAT_OUT, O 
                           => G_3215GAT_OUT);
   G_3212GAT : Nor_gate port map( I1 => G_3145GAT_OUT, I2 => G_3146GAT_OUT, O 
                           => G_3212GAT_OUT);
   G_3208GAT : Nor_gate port map( I1 => G_2983GAT_OUT, I2 => G_3136GAT_OUT, O 
                           => G_3208GAT_OUT);
   G_3207GAT : Nor_gate port map( I1 => G_3136GAT_OUT, I2 => G_1236GAT_OUT, O 
                           => G_3207GAT_OUT);
   G_3206GAT : Nor_gate port map( I1 => G_3076GAT_OUT, I2 => G_3136GAT_OUT, O 
                           => G_3206GAT_OUT);
   G_3202GAT : Nor_gate port map( I1 => G_3133GAT_OUT, I2 => G_1188GAT_OUT, O 
                           => G_3202GAT_OUT);
   G_3199GAT : Nor_gate port map( I1 => G_3131GAT_OUT, I2 => G_3132GAT_OUT, O 
                           => G_3199GAT_OUT);
   G_3198GAT : Nor_gate port map( I1 => G_3127GAT_OUT, I2 => G_3064GAT_OUT, O 
                           => G_3198GAT_OUT);
   G_3197GAT : Nor_gate port map( I1 => G_3067GAT_OUT, I2 => G_3127GAT_OUT, O 
                           => G_3197GAT_OUT);
   G_3193GAT : Nor_gate port map( I1 => G_3124GAT_OUT, I2 => G_3121GAT_OUT, O 
                           => G_3193GAT_OUT);
   G_3190GAT : Nor_gate port map( I1 => G_3119GAT_OUT, I2 => G_3120GAT_OUT, O 
                           => G_3190GAT_OUT);
   G_3187GAT : Nor_gate port map( I1 => G_2962GAT_OUT, I2 => G_3115GAT_OUT, O 
                           => G_3187GAT_OUT);
   G_3186GAT : Nor_gate port map( I1 => G_3115GAT_OUT, I2 => G_993GAT_OUT, O =>
                           G_3186GAT_OUT);
   G_3185GAT : Nor_gate port map( I1 => G_3055GAT_OUT, I2 => G_3115GAT_OUT, O 
                           => G_3185GAT_OUT);
   G_3182GAT : Nor_gate port map( I1 => G_2958GAT_OUT, I2 => G_3111GAT_OUT, O 
                           => G_3182GAT_OUT);
   G_3181GAT : Nor_gate port map( I1 => G_3111GAT_OUT, I2 => G_945GAT_OUT, O =>
                           G_3181GAT_OUT);
   G_3180GAT : Nor_gate port map( I1 => G_3052GAT_OUT, I2 => G_3111GAT_OUT, O 
                           => G_3180GAT_OUT);
   G_3177GAT : Nor_gate port map( I1 => G_2954GAT_OUT, I2 => G_3107GAT_OUT, O 
                           => G_3177GAT_OUT);
   G_3176GAT : Nor_gate port map( I1 => G_3107GAT_OUT, I2 => G_897GAT_OUT, O =>
                           G_3176GAT_OUT);
   G_3175GAT : Nor_gate port map( I1 => G_3049GAT_OUT, I2 => G_3107GAT_OUT, O 
                           => G_3175GAT_OUT);
   G_3172GAT : Nor_gate port map( I1 => G_2950GAT_OUT, I2 => G_3103GAT_OUT, O 
                           => G_3172GAT_OUT);
   G_3171GAT : Nor_gate port map( I1 => G_3103GAT_OUT, I2 => G_849GAT_OUT, O =>
                           G_3171GAT_OUT);
   G_3170GAT : Nor_gate port map( I1 => G_3046GAT_OUT, I2 => G_3103GAT_OUT, O 
                           => G_3170GAT_OUT);
   G_3167GAT : Nor_gate port map( I1 => G_2946GAT_OUT, I2 => G_3099GAT_OUT, O 
                           => G_3167GAT_OUT);
   G_3166GAT : Nor_gate port map( I1 => G_3099GAT_OUT, I2 => G_801GAT_OUT, O =>
                           G_3166GAT_OUT);
   G_3165GAT : Nor_gate port map( I1 => G_3043GAT_OUT, I2 => G_3099GAT_OUT, O 
                           => G_3165GAT_OUT);
   G_3162GAT : Nor_gate port map( I1 => G_2942GAT_OUT, I2 => G_3095GAT_OUT, O 
                           => G_3162GAT_OUT);
   G_3161GAT : Nor_gate port map( I1 => G_3095GAT_OUT, I2 => G_753GAT_OUT, O =>
                           G_3161GAT_OUT);
   G_3160GAT : Nor_gate port map( I1 => G_3040GAT_OUT, I2 => G_3095GAT_OUT, O 
                           => G_3160GAT_OUT);
   G_3157GAT : Nor_gate port map( I1 => G_2938GAT_OUT, I2 => G_3091GAT_OUT, O 
                           => G_3157GAT_OUT);
   G_3156GAT : Nor_gate port map( I1 => G_3091GAT_OUT, I2 => G_705GAT_OUT, O =>
                           G_3156GAT_OUT);
   G_3155GAT : Nor_gate port map( I1 => G_3037GAT_OUT, I2 => G_3091GAT_OUT, O 
                           => G_3155GAT_OUT);
   G_3152GAT : Nor_gate port map( I1 => G_2934GAT_OUT, I2 => G_3087GAT_OUT, O 
                           => G_3152GAT_OUT);
   G_3151GAT : Nor_gate port map( I1 => G_3087GAT_OUT, I2 => G_657GAT_OUT, O =>
                           G_3151GAT_OUT);
   G_3150GAT : Nor_gate port map( I1 => G_3034GAT_OUT, I2 => G_3087GAT_OUT, O 
                           => G_3150GAT_OUT);
   G_3147GAT : Nor_gate port map( I1 => G_2930GAT_OUT, I2 => G_3083GAT_OUT, O 
                           => G_3147GAT_OUT);
   G_3146GAT : Nor_gate port map( I1 => G_3083GAT_OUT, I2 => G_609GAT_OUT, O =>
                           G_3146GAT_OUT);
   G_3145GAT : Nor_gate port map( I1 => G_3031GAT_OUT, I2 => G_3083GAT_OUT, O 
                           => G_3145GAT_OUT);
   G_3142GAT : Nor_gate port map( I1 => G_2926GAT_OUT, I2 => G_3079GAT_OUT, O 
                           => G_3142GAT_OUT);
   G_3141GAT : Nor_gate port map( I1 => G_3079GAT_OUT, I2 => G_561GAT_OUT, O =>
                           G_3141GAT_OUT);
   G_3140GAT : Nor_gate port map( I1 => G_3028GAT_OUT, I2 => G_3079GAT_OUT, O 
                           => G_3140GAT_OUT);
   G_3136GAT : Nor_gate port map( I1 => G_3076GAT_OUT, I2 => G_1236GAT_OUT, O 
                           => G_3136GAT_OUT);
   G_3133GAT : Nor_gate port map( I1 => G_3074GAT_OUT, I2 => G_3075GAT_OUT, O 
                           => G_3133GAT_OUT);
   G_3132GAT : Nor_gate port map( I1 => G_3070GAT_OUT, I2 => G_3016GAT_OUT, O 
                           => G_3132GAT_OUT);
   G_3131GAT : Nor_gate port map( I1 => G_3019GAT_OUT, I2 => G_3070GAT_OUT, O 
                           => G_3131GAT_OUT);
   G_3127GAT : Nor_gate port map( I1 => G_3067GAT_OUT, I2 => G_3064GAT_OUT, O 
                           => G_3127GAT_OUT);
   G_3124GAT : Nor_gate port map( I1 => G_3062GAT_OUT, I2 => G_3063GAT_OUT, O 
                           => G_3124GAT_OUT);
   G_3121GAT : Nor_gate port map( I1 => G_2908GAT_OUT, I2 => G_3058GAT_OUT, O 
                           => G_3121GAT_OUT);
   G_3120GAT : Nor_gate port map( I1 => G_3058GAT_OUT, I2 => G_1041GAT_OUT, O 
                           => G_3120GAT_OUT);
   G_3119GAT : Nor_gate port map( I1 => G_3007GAT_OUT, I2 => G_3058GAT_OUT, O 
                           => G_3119GAT_OUT);
   G_3115GAT : Nor_gate port map( I1 => G_3055GAT_OUT, I2 => G_993GAT_OUT, O =>
                           G_3115GAT_OUT);
   G_3111GAT : Nor_gate port map( I1 => G_3052GAT_OUT, I2 => G_945GAT_OUT, O =>
                           G_3111GAT_OUT);
   G_3107GAT : Nor_gate port map( I1 => G_3049GAT_OUT, I2 => G_897GAT_OUT, O =>
                           G_3107GAT_OUT);
   G_3103GAT : Nor_gate port map( I1 => G_3046GAT_OUT, I2 => G_849GAT_OUT, O =>
                           G_3103GAT_OUT);
   G_3099GAT : Nor_gate port map( I1 => G_3043GAT_OUT, I2 => G_801GAT_OUT, O =>
                           G_3099GAT_OUT);
   G_3095GAT : Nor_gate port map( I1 => G_3040GAT_OUT, I2 => G_753GAT_OUT, O =>
                           G_3095GAT_OUT);
   G_3091GAT : Nor_gate port map( I1 => G_3037GAT_OUT, I2 => G_705GAT_OUT, O =>
                           G_3091GAT_OUT);
   G_3087GAT : Nor_gate port map( I1 => G_3034GAT_OUT, I2 => G_657GAT_OUT, O =>
                           G_3087GAT_OUT);
   G_3083GAT : Nor_gate port map( I1 => G_3031GAT_OUT, I2 => G_609GAT_OUT, O =>
                           G_3083GAT_OUT);
   G_3079GAT : Nor_gate port map( I1 => G_3028GAT_OUT, I2 => G_561GAT_OUT, O =>
                           G_3079GAT_OUT);
   G_3076GAT : Nor_gate port map( I1 => G_3026GAT_OUT, I2 => G_3027GAT_OUT, O 
                           => G_3076GAT_OUT);
   G_3075GAT : Nor_gate port map( I1 => G_3022GAT_OUT, I2 => G_2977GAT_OUT, O 
                           => G_3075GAT_OUT);
   G_3074GAT : Nor_gate port map( I1 => G_2980GAT_OUT, I2 => G_3022GAT_OUT, O 
                           => G_3074GAT_OUT);
   G_3070GAT : Nor_gate port map( I1 => G_3019GAT_OUT, I2 => G_3016GAT_OUT, O 
                           => G_3070GAT_OUT);
   G_3067GAT : Nor_gate port map( I1 => G_3014GAT_OUT, I2 => G_3015GAT_OUT, O 
                           => G_3067GAT_OUT);
   G_3064GAT : Nor_gate port map( I1 => G_2864GAT_OUT, I2 => G_3010GAT_OUT, O 
                           => G_3064GAT_OUT);
   G_3063GAT : Nor_gate port map( I1 => G_3010GAT_OUT, I2 => G_1089GAT_OUT, O 
                           => G_3063GAT_OUT);
   G_3062GAT : Nor_gate port map( I1 => G_2968GAT_OUT, I2 => G_3010GAT_OUT, O 
                           => G_3062GAT_OUT);
   G_3058GAT : Nor_gate port map( I1 => G_3007GAT_OUT, I2 => G_1041GAT_OUT, O 
                           => G_3058GAT_OUT);
   G_3055GAT : Nor_gate port map( I1 => G_3005GAT_OUT, I2 => G_3006GAT_OUT, O 
                           => G_3055GAT_OUT);
   G_3052GAT : Nor_gate port map( I1 => G_3003GAT_OUT, I2 => G_3004GAT_OUT, O 
                           => G_3052GAT_OUT);
   G_3049GAT : Nor_gate port map( I1 => G_3001GAT_OUT, I2 => G_3002GAT_OUT, O 
                           => G_3049GAT_OUT);
   G_3046GAT : Nor_gate port map( I1 => G_2999GAT_OUT, I2 => G_3000GAT_OUT, O 
                           => G_3046GAT_OUT);
   G_3043GAT : Nor_gate port map( I1 => G_2997GAT_OUT, I2 => G_2998GAT_OUT, O 
                           => G_3043GAT_OUT);
   G_3040GAT : Nor_gate port map( I1 => G_2995GAT_OUT, I2 => G_2996GAT_OUT, O 
                           => G_3040GAT_OUT);
   G_3037GAT : Nor_gate port map( I1 => G_2993GAT_OUT, I2 => G_2994GAT_OUT, O 
                           => G_3037GAT_OUT);
   G_3034GAT : Nor_gate port map( I1 => G_2991GAT_OUT, I2 => G_2992GAT_OUT, O 
                           => G_3034GAT_OUT);
   G_3031GAT : Nor_gate port map( I1 => G_2989GAT_OUT, I2 => G_2990GAT_OUT, O 
                           => G_3031GAT_OUT);
   G_3028GAT : Nor_gate port map( I1 => G_2987GAT_OUT, I2 => G_2988GAT_OUT, O 
                           => G_3028GAT_OUT);
   G_3027GAT : Nor_gate port map( I1 => G_2983GAT_OUT, I2 => G_2923GAT_OUT, O 
                           => G_3027GAT_OUT);
   G_3026GAT : Nor_gate port map( I1 => G_1281GAT_OUT, I2 => G_2983GAT_OUT, O 
                           => G_3026GAT_OUT);
   G_3022GAT : Nor_gate port map( I1 => G_2980GAT_OUT, I2 => G_2977GAT_OUT, O 
                           => G_3022GAT_OUT);
   G_3019GAT : Nor_gate port map( I1 => G_2975GAT_OUT, I2 => G_2976GAT_OUT, O 
                           => G_3019GAT_OUT);
   G_3016GAT : Nor_gate port map( I1 => G_2797GAT_OUT, I2 => G_2971GAT_OUT, O 
                           => G_3016GAT_OUT);
   G_3015GAT : Nor_gate port map( I1 => G_2971GAT_OUT, I2 => G_1137GAT_OUT, O 
                           => G_3015GAT_OUT);
   G_3014GAT : Nor_gate port map( I1 => G_2914GAT_OUT, I2 => G_2971GAT_OUT, O 
                           => G_3014GAT_OUT);
   G_3010GAT : Nor_gate port map( I1 => G_2968GAT_OUT, I2 => G_1089GAT_OUT, O 
                           => G_3010GAT_OUT);
   G_3007GAT : Nor_gate port map( I1 => G_2966GAT_OUT, I2 => G_2967GAT_OUT, O 
                           => G_3007GAT_OUT);
   G_3006GAT : Nor_gate port map( I1 => G_2962GAT_OUT, I2 => G_2853GAT_OUT, O 
                           => G_3006GAT_OUT);
   G_3005GAT : Nor_gate port map( I1 => G_2905GAT_OUT, I2 => G_2962GAT_OUT, O 
                           => G_3005GAT_OUT);
   G_3004GAT : Nor_gate port map( I1 => G_2958GAT_OUT, I2 => G_2848GAT_OUT, O 
                           => G_3004GAT_OUT);
   G_3003GAT : Nor_gate port map( I1 => G_2902GAT_OUT, I2 => G_2958GAT_OUT, O 
                           => G_3003GAT_OUT);
   G_3002GAT : Nor_gate port map( I1 => G_2954GAT_OUT, I2 => G_2843GAT_OUT, O 
                           => G_3002GAT_OUT);
   G_3001GAT : Nor_gate port map( I1 => G_2899GAT_OUT, I2 => G_2954GAT_OUT, O 
                           => G_3001GAT_OUT);
   G_3000GAT : Nor_gate port map( I1 => G_2950GAT_OUT, I2 => G_2838GAT_OUT, O 
                           => G_3000GAT_OUT);
   G_2999GAT : Nor_gate port map( I1 => G_2896GAT_OUT, I2 => G_2950GAT_OUT, O 
                           => G_2999GAT_OUT);
   G_2998GAT : Nor_gate port map( I1 => G_2946GAT_OUT, I2 => G_2833GAT_OUT, O 
                           => G_2998GAT_OUT);
   G_2997GAT : Nor_gate port map( I1 => G_2893GAT_OUT, I2 => G_2946GAT_OUT, O 
                           => G_2997GAT_OUT);
   G_2996GAT : Nor_gate port map( I1 => G_2942GAT_OUT, I2 => G_2828GAT_OUT, O 
                           => G_2996GAT_OUT);
   G_2995GAT : Nor_gate port map( I1 => G_2890GAT_OUT, I2 => G_2942GAT_OUT, O 
                           => G_2995GAT_OUT);
   G_2994GAT : Nor_gate port map( I1 => G_2938GAT_OUT, I2 => G_2823GAT_OUT, O 
                           => G_2994GAT_OUT);
   G_2993GAT : Nor_gate port map( I1 => G_2887GAT_OUT, I2 => G_2938GAT_OUT, O 
                           => G_2993GAT_OUT);
   G_2992GAT : Nor_gate port map( I1 => G_2934GAT_OUT, I2 => G_2818GAT_OUT, O 
                           => G_2992GAT_OUT);
   G_2991GAT : Nor_gate port map( I1 => G_2884GAT_OUT, I2 => G_2934GAT_OUT, O 
                           => G_2991GAT_OUT);
   G_2990GAT : Nor_gate port map( I1 => G_2930GAT_OUT, I2 => G_2813GAT_OUT, O 
                           => G_2990GAT_OUT);
   G_2989GAT : Nor_gate port map( I1 => G_2881GAT_OUT, I2 => G_2930GAT_OUT, O 
                           => G_2989GAT_OUT);
   G_2988GAT : Nor_gate port map( I1 => G_2926GAT_OUT, I2 => G_2808GAT_OUT, O 
                           => G_2988GAT_OUT);
   G_2987GAT : Nor_gate port map( I1 => G_2878GAT_OUT, I2 => G_2926GAT_OUT, O 
                           => G_2987GAT_OUT);
   G_2983GAT : Nor_gate port map( I1 => G_1281GAT_OUT, I2 => G_2923GAT_OUT, O 
                           => G_2983GAT_OUT);
   G_2980GAT : Nor_gate port map( I1 => G_2921GAT_OUT, I2 => G_2922GAT_OUT, O 
                           => G_2980GAT_OUT);
   G_2977GAT : Nor_gate port map( I1 => G_2739GAT_OUT, I2 => G_2917GAT_OUT, O 
                           => G_2977GAT_OUT);
   G_2976GAT : Nor_gate port map( I1 => G_2917GAT_OUT, I2 => G_1185GAT_OUT, O 
                           => G_2976GAT_OUT);
   G_2975GAT : Nor_gate port map( I1 => G_2870GAT_OUT, I2 => G_2917GAT_OUT, O 
                           => G_2975GAT_OUT);
   G_2971GAT : Nor_gate port map( I1 => G_2914GAT_OUT, I2 => G_1137GAT_OUT, O 
                           => G_2971GAT_OUT);
   G_2968GAT : Nor_gate port map( I1 => G_2912GAT_OUT, I2 => G_2913GAT_OUT, O 
                           => G_2968GAT_OUT);
   G_2967GAT : Nor_gate port map( I1 => G_2908GAT_OUT, I2 => G_2858GAT_OUT, O 
                           => G_2967GAT_OUT);
   G_2966GAT : Nor_gate port map( I1 => G_2861GAT_OUT, I2 => G_2908GAT_OUT, O 
                           => G_2966GAT_OUT);
   G_2962GAT : Nor_gate port map( I1 => G_2905GAT_OUT, I2 => G_2853GAT_OUT, O 
                           => G_2962GAT_OUT);
   G_2958GAT : Nor_gate port map( I1 => G_2902GAT_OUT, I2 => G_2848GAT_OUT, O 
                           => G_2958GAT_OUT);
   G_2954GAT : Nor_gate port map( I1 => G_2899GAT_OUT, I2 => G_2843GAT_OUT, O 
                           => G_2954GAT_OUT);
   G_2950GAT : Nor_gate port map( I1 => G_2896GAT_OUT, I2 => G_2838GAT_OUT, O 
                           => G_2950GAT_OUT);
   G_2946GAT : Nor_gate port map( I1 => G_2893GAT_OUT, I2 => G_2833GAT_OUT, O 
                           => G_2946GAT_OUT);
   G_2942GAT : Nor_gate port map( I1 => G_2890GAT_OUT, I2 => G_2828GAT_OUT, O 
                           => G_2942GAT_OUT);
   G_2938GAT : Nor_gate port map( I1 => G_2887GAT_OUT, I2 => G_2823GAT_OUT, O 
                           => G_2938GAT_OUT);
   G_2934GAT : Nor_gate port map( I1 => G_2884GAT_OUT, I2 => G_2818GAT_OUT, O 
                           => G_2934GAT_OUT);
   G_2930GAT : Nor_gate port map( I1 => G_2881GAT_OUT, I2 => G_2813GAT_OUT, O 
                           => G_2930GAT_OUT);
   G_2926GAT : Nor_gate port map( I1 => G_2878GAT_OUT, I2 => G_2808GAT_OUT, O 
                           => G_2926GAT_OUT);
   G_2923GAT : Nor_gate port map( I1 => G_2690GAT_OUT, I2 => G_2873GAT_OUT, O 
                           => G_2923GAT_OUT);
   G_2922GAT : Nor_gate port map( I1 => G_2873GAT_OUT, I2 => G_1233GAT_OUT, O 
                           => G_2922GAT_OUT);
   G_2921GAT : Nor_gate port map( I1 => G_2803GAT_OUT, I2 => G_2873GAT_OUT, O 
                           => G_2921GAT_OUT);
   G_2917GAT : Nor_gate port map( I1 => G_2870GAT_OUT, I2 => G_1185GAT_OUT, O 
                           => G_2917GAT_OUT);
   G_2914GAT : Nor_gate port map( I1 => G_2868GAT_OUT, I2 => G_2869GAT_OUT, O 
                           => G_2914GAT_OUT);
   G_2913GAT : Nor_gate port map( I1 => G_2864GAT_OUT, I2 => G_2791GAT_OUT, O 
                           => G_2913GAT_OUT);
   G_2912GAT : Nor_gate port map( I1 => G_2794GAT_OUT, I2 => G_2864GAT_OUT, O 
                           => G_2912GAT_OUT);
   G_2908GAT : Nor_gate port map( I1 => G_2861GAT_OUT, I2 => G_2858GAT_OUT, O 
                           => G_2908GAT_OUT);
   G_2905GAT : Nor_gate port map( I1 => G_2856GAT_OUT, I2 => G_2857GAT_OUT, O 
                           => G_2905GAT_OUT);
   G_2902GAT : Nor_gate port map( I1 => G_2851GAT_OUT, I2 => G_2852GAT_OUT, O 
                           => G_2902GAT_OUT);
   G_2899GAT : Nor_gate port map( I1 => G_2846GAT_OUT, I2 => G_2847GAT_OUT, O 
                           => G_2899GAT_OUT);
   G_2896GAT : Nor_gate port map( I1 => G_2841GAT_OUT, I2 => G_2842GAT_OUT, O 
                           => G_2896GAT_OUT);
   G_2893GAT : Nor_gate port map( I1 => G_2836GAT_OUT, I2 => G_2837GAT_OUT, O 
                           => G_2893GAT_OUT);
   G_2890GAT : Nor_gate port map( I1 => G_2831GAT_OUT, I2 => G_2832GAT_OUT, O 
                           => G_2890GAT_OUT);
   G_2887GAT : Nor_gate port map( I1 => G_2826GAT_OUT, I2 => G_2827GAT_OUT, O 
                           => G_2887GAT_OUT);
   G_2884GAT : Nor_gate port map( I1 => G_2821GAT_OUT, I2 => G_2822GAT_OUT, O 
                           => G_2884GAT_OUT);
   G_2881GAT : Nor_gate port map( I1 => G_2816GAT_OUT, I2 => G_2817GAT_OUT, O 
                           => G_2881GAT_OUT);
   G_2878GAT : Nor_gate port map( I1 => G_2811GAT_OUT, I2 => G_2812GAT_OUT, O 
                           => G_2878GAT_OUT);
   G_2873GAT : Nor_gate port map( I1 => G_2803GAT_OUT, I2 => G_1233GAT_OUT, O 
                           => G_2873GAT_OUT);
   G_2870GAT : Nor_gate port map( I1 => G_2801GAT_OUT, I2 => G_2802GAT_OUT, O 
                           => G_2870GAT_OUT);
   G_2869GAT : Nor_gate port map( I1 => G_2797GAT_OUT, I2 => G_2733GAT_OUT, O 
                           => G_2869GAT_OUT);
   G_2868GAT : Nor_gate port map( I1 => G_2736GAT_OUT, I2 => G_2797GAT_OUT, O 
                           => G_2868GAT_OUT);
   G_2864GAT : Nor_gate port map( I1 => G_2794GAT_OUT, I2 => G_2791GAT_OUT, O 
                           => G_2864GAT_OUT);
   G_2861GAT : Nor_gate port map( I1 => G_2789GAT_OUT, I2 => G_2790GAT_OUT, O 
                           => G_2861GAT_OUT);
   G_2858GAT : Nor_gate port map( I1 => G_2635GAT_OUT, I2 => G_2785GAT_OUT, O 
                           => G_2858GAT_OUT);
   G_2857GAT : Nor_gate port map( I1 => G_2785GAT_OUT, I2 => G_1038GAT_OUT, O 
                           => G_2857GAT_OUT);
   G_2856GAT : Nor_gate port map( I1 => G_2724GAT_OUT, I2 => G_2785GAT_OUT, O 
                           => G_2856GAT_OUT);
   G_2853GAT : Nor_gate port map( I1 => G_2631GAT_OUT, I2 => G_2781GAT_OUT, O 
                           => G_2853GAT_OUT);
   G_2852GAT : Nor_gate port map( I1 => G_2781GAT_OUT, I2 => G_990GAT_OUT, O =>
                           G_2852GAT_OUT);
   G_2851GAT : Nor_gate port map( I1 => G_2721GAT_OUT, I2 => G_2781GAT_OUT, O 
                           => G_2851GAT_OUT);
   G_2848GAT : Nor_gate port map( I1 => G_2627GAT_OUT, I2 => G_2777GAT_OUT, O 
                           => G_2848GAT_OUT);
   G_2847GAT : Nor_gate port map( I1 => G_2777GAT_OUT, I2 => G_942GAT_OUT, O =>
                           G_2847GAT_OUT);
   G_2846GAT : Nor_gate port map( I1 => G_2718GAT_OUT, I2 => G_2777GAT_OUT, O 
                           => G_2846GAT_OUT);
   G_2843GAT : Nor_gate port map( I1 => G_2623GAT_OUT, I2 => G_2773GAT_OUT, O 
                           => G_2843GAT_OUT);
   G_2842GAT : Nor_gate port map( I1 => G_2773GAT_OUT, I2 => G_894GAT_OUT, O =>
                           G_2842GAT_OUT);
   G_2841GAT : Nor_gate port map( I1 => G_2715GAT_OUT, I2 => G_2773GAT_OUT, O 
                           => G_2841GAT_OUT);
   G_2838GAT : Nor_gate port map( I1 => G_2619GAT_OUT, I2 => G_2769GAT_OUT, O 
                           => G_2838GAT_OUT);
   G_2837GAT : Nor_gate port map( I1 => G_2769GAT_OUT, I2 => G_846GAT_OUT, O =>
                           G_2837GAT_OUT);
   G_2836GAT : Nor_gate port map( I1 => G_2712GAT_OUT, I2 => G_2769GAT_OUT, O 
                           => G_2836GAT_OUT);
   G_2833GAT : Nor_gate port map( I1 => G_2615GAT_OUT, I2 => G_2765GAT_OUT, O 
                           => G_2833GAT_OUT);
   G_2832GAT : Nor_gate port map( I1 => G_2765GAT_OUT, I2 => G_798GAT_OUT, O =>
                           G_2832GAT_OUT);
   G_2831GAT : Nor_gate port map( I1 => G_2709GAT_OUT, I2 => G_2765GAT_OUT, O 
                           => G_2831GAT_OUT);
   G_2828GAT : Nor_gate port map( I1 => G_2611GAT_OUT, I2 => G_2761GAT_OUT, O 
                           => G_2828GAT_OUT);
   G_2827GAT : Nor_gate port map( I1 => G_2761GAT_OUT, I2 => G_750GAT_OUT, O =>
                           G_2827GAT_OUT);
   G_2826GAT : Nor_gate port map( I1 => G_2706GAT_OUT, I2 => G_2761GAT_OUT, O 
                           => G_2826GAT_OUT);
   G_2823GAT : Nor_gate port map( I1 => G_2607GAT_OUT, I2 => G_2757GAT_OUT, O 
                           => G_2823GAT_OUT);
   G_2822GAT : Nor_gate port map( I1 => G_2757GAT_OUT, I2 => G_702GAT_OUT, O =>
                           G_2822GAT_OUT);
   G_2821GAT : Nor_gate port map( I1 => G_2703GAT_OUT, I2 => G_2757GAT_OUT, O 
                           => G_2821GAT_OUT);
   G_2818GAT : Nor_gate port map( I1 => G_2603GAT_OUT, I2 => G_2753GAT_OUT, O 
                           => G_2818GAT_OUT);
   G_2817GAT : Nor_gate port map( I1 => G_2753GAT_OUT, I2 => G_654GAT_OUT, O =>
                           G_2817GAT_OUT);
   G_2816GAT : Nor_gate port map( I1 => G_2700GAT_OUT, I2 => G_2753GAT_OUT, O 
                           => G_2816GAT_OUT);
   G_2813GAT : Nor_gate port map( I1 => G_2599GAT_OUT, I2 => G_2749GAT_OUT, O 
                           => G_2813GAT_OUT);
   G_2812GAT : Nor_gate port map( I1 => G_2749GAT_OUT, I2 => G_606GAT_OUT, O =>
                           G_2812GAT_OUT);
   G_2811GAT : Nor_gate port map( I1 => G_2697GAT_OUT, I2 => G_2749GAT_OUT, O 
                           => G_2811GAT_OUT);
   G_2808GAT : Nor_gate port map( I1 => G_2595GAT_OUT, I2 => G_2745GAT_OUT, O 
                           => G_2808GAT_OUT);
   G_2807GAT : Nor_gate port map( I1 => G_2745GAT_OUT, I2 => G_558GAT_OUT, O =>
                           G_2807GAT_OUT);
   G_2806GAT : Nor_gate port map( I1 => G_2694GAT_OUT, I2 => G_2745GAT_OUT, O 
                           => G_2806GAT_OUT);
   G_2803GAT : Nor_gate port map( I1 => G_2743GAT_OUT, I2 => G_2744GAT_OUT, O 
                           => G_2803GAT_OUT);
   G_2802GAT : Nor_gate port map( I1 => G_2739GAT_OUT, I2 => G_2684GAT_OUT, O 
                           => G_2802GAT_OUT);
   G_2801GAT : Nor_gate port map( I1 => G_2687GAT_OUT, I2 => G_2739GAT_OUT, O 
                           => G_2801GAT_OUT);
   G_2797GAT : Nor_gate port map( I1 => G_2736GAT_OUT, I2 => G_2733GAT_OUT, O 
                           => G_2797GAT_OUT);
   G_2794GAT : Nor_gate port map( I1 => G_2731GAT_OUT, I2 => G_2732GAT_OUT, O 
                           => G_2794GAT_OUT);
   G_2791GAT : Nor_gate port map( I1 => G_2582GAT_OUT, I2 => G_2727GAT_OUT, O 
                           => G_2791GAT_OUT);
   G_2790GAT : Nor_gate port map( I1 => G_2727GAT_OUT, I2 => G_1086GAT_OUT, O 
                           => G_2790GAT_OUT);
   G_2789GAT : Nor_gate port map( I1 => G_2675GAT_OUT, I2 => G_2727GAT_OUT, O 
                           => G_2789GAT_OUT);
   G_2785GAT : Nor_gate port map( I1 => G_2724GAT_OUT, I2 => G_1038GAT_OUT, O 
                           => G_2785GAT_OUT);
   G_2781GAT : Nor_gate port map( I1 => G_2721GAT_OUT, I2 => G_990GAT_OUT, O =>
                           G_2781GAT_OUT);
   G_2777GAT : Nor_gate port map( I1 => G_2718GAT_OUT, I2 => G_942GAT_OUT, O =>
                           G_2777GAT_OUT);
   G_2773GAT : Nor_gate port map( I1 => G_2715GAT_OUT, I2 => G_894GAT_OUT, O =>
                           G_2773GAT_OUT);
   G_2769GAT : Nor_gate port map( I1 => G_2712GAT_OUT, I2 => G_846GAT_OUT, O =>
                           G_2769GAT_OUT);
   G_2765GAT : Nor_gate port map( I1 => G_2709GAT_OUT, I2 => G_798GAT_OUT, O =>
                           G_2765GAT_OUT);
   G_2761GAT : Nor_gate port map( I1 => G_2706GAT_OUT, I2 => G_750GAT_OUT, O =>
                           G_2761GAT_OUT);
   G_2757GAT : Nor_gate port map( I1 => G_2703GAT_OUT, I2 => G_702GAT_OUT, O =>
                           G_2757GAT_OUT);
   G_2753GAT : Nor_gate port map( I1 => G_2700GAT_OUT, I2 => G_654GAT_OUT, O =>
                           G_2753GAT_OUT);
   G_2749GAT : Nor_gate port map( I1 => G_2697GAT_OUT, I2 => G_606GAT_OUT, O =>
                           G_2749GAT_OUT);
   G_2745GAT : Nor_gate port map( I1 => G_2694GAT_OUT, I2 => G_558GAT_OUT, O =>
                           G_2745GAT_OUT);
   G_2744GAT : Nor_gate port map( I1 => G_2690GAT_OUT, I2 => G_2650GAT_OUT, O 
                           => G_2744GAT_OUT);
   G_2743GAT : Nor_gate port map( I1 => G_1278GAT_OUT, I2 => G_2690GAT_OUT, O 
                           => G_2743GAT_OUT);
   G_2739GAT : Nor_gate port map( I1 => G_2687GAT_OUT, I2 => G_2684GAT_OUT, O 
                           => G_2739GAT_OUT);
   G_2736GAT : Nor_gate port map( I1 => G_2682GAT_OUT, I2 => G_2683GAT_OUT, O 
                           => G_2736GAT_OUT);
   G_2733GAT : Nor_gate port map( I1 => G_2539GAT_OUT, I2 => G_2678GAT_OUT, O 
                           => G_2733GAT_OUT);
   G_2732GAT : Nor_gate port map( I1 => G_2678GAT_OUT, I2 => G_1134GAT_OUT, O 
                           => G_2732GAT_OUT);
   G_2731GAT : Nor_gate port map( I1 => G_2641GAT_OUT, I2 => G_2678GAT_OUT, O 
                           => G_2731GAT_OUT);
   G_2727GAT : Nor_gate port map( I1 => G_2675GAT_OUT, I2 => G_1086GAT_OUT, O 
                           => G_2727GAT_OUT);
   G_2724GAT : Nor_gate port map( I1 => G_2673GAT_OUT, I2 => G_2674GAT_OUT, O 
                           => G_2724GAT_OUT);
   G_2721GAT : Nor_gate port map( I1 => G_2671GAT_OUT, I2 => G_2672GAT_OUT, O 
                           => G_2721GAT_OUT);
   G_2718GAT : Nor_gate port map( I1 => G_2669GAT_OUT, I2 => G_2670GAT_OUT, O 
                           => G_2718GAT_OUT);
   G_2715GAT : Nor_gate port map( I1 => G_2667GAT_OUT, I2 => G_2668GAT_OUT, O 
                           => G_2715GAT_OUT);
   G_2712GAT : Nor_gate port map( I1 => G_2665GAT_OUT, I2 => G_2666GAT_OUT, O 
                           => G_2712GAT_OUT);
   G_2709GAT : Nor_gate port map( I1 => G_2663GAT_OUT, I2 => G_2664GAT_OUT, O 
                           => G_2709GAT_OUT);
   G_2706GAT : Nor_gate port map( I1 => G_2661GAT_OUT, I2 => G_2662GAT_OUT, O 
                           => G_2706GAT_OUT);
   G_2703GAT : Nor_gate port map( I1 => G_2659GAT_OUT, I2 => G_2660GAT_OUT, O 
                           => G_2703GAT_OUT);
   G_2700GAT : Nor_gate port map( I1 => G_2657GAT_OUT, I2 => G_2658GAT_OUT, O 
                           => G_2700GAT_OUT);
   G_2697GAT : Nor_gate port map( I1 => G_2655GAT_OUT, I2 => G_2656GAT_OUT, O 
                           => G_2697GAT_OUT);
   G_2694GAT : Nor_gate port map( I1 => G_2653GAT_OUT, I2 => G_2654GAT_OUT, O 
                           => G_2694GAT_OUT);
   G_2690GAT : Nor_gate port map( I1 => G_1278GAT_OUT, I2 => G_2650GAT_OUT, O 
                           => G_2690GAT_OUT);
   G_2687GAT : Nor_gate port map( I1 => G_2648GAT_OUT, I2 => G_2649GAT_OUT, O 
                           => G_2687GAT_OUT);
   G_2684GAT : Nor_gate port map( I1 => G_2470GAT_OUT, I2 => G_2644GAT_OUT, O 
                           => G_2684GAT_OUT);
   G_2683GAT : Nor_gate port map( I1 => G_2644GAT_OUT, I2 => G_1182GAT_OUT, O 
                           => G_2683GAT_OUT);
   G_2682GAT : Nor_gate port map( I1 => G_2588GAT_OUT, I2 => G_2644GAT_OUT, O 
                           => G_2682GAT_OUT);
   G_2678GAT : Nor_gate port map( I1 => G_2641GAT_OUT, I2 => G_1134GAT_OUT, O 
                           => G_2678GAT_OUT);
   G_2675GAT : Nor_gate port map( I1 => G_2639GAT_OUT, I2 => G_2640GAT_OUT, O 
                           => G_2675GAT_OUT);
   G_2674GAT : Nor_gate port map( I1 => G_2635GAT_OUT, I2 => G_2528GAT_OUT, O 
                           => G_2674GAT_OUT);
   G_2673GAT : Nor_gate port map( I1 => G_2579GAT_OUT, I2 => G_2635GAT_OUT, O 
                           => G_2673GAT_OUT);
   G_2672GAT : Nor_gate port map( I1 => G_2631GAT_OUT, I2 => G_2523GAT_OUT, O 
                           => G_2672GAT_OUT);
   G_2671GAT : Nor_gate port map( I1 => G_2576GAT_OUT, I2 => G_2631GAT_OUT, O 
                           => G_2671GAT_OUT);
   G_2670GAT : Nor_gate port map( I1 => G_2627GAT_OUT, I2 => G_2518GAT_OUT, O 
                           => G_2670GAT_OUT);
   G_2669GAT : Nor_gate port map( I1 => G_2573GAT_OUT, I2 => G_2627GAT_OUT, O 
                           => G_2669GAT_OUT);
   G_2668GAT : Nor_gate port map( I1 => G_2623GAT_OUT, I2 => G_2513GAT_OUT, O 
                           => G_2668GAT_OUT);
   G_2667GAT : Nor_gate port map( I1 => G_2570GAT_OUT, I2 => G_2623GAT_OUT, O 
                           => G_2667GAT_OUT);
   G_2666GAT : Nor_gate port map( I1 => G_2619GAT_OUT, I2 => G_2508GAT_OUT, O 
                           => G_2666GAT_OUT);
   G_2665GAT : Nor_gate port map( I1 => G_2567GAT_OUT, I2 => G_2619GAT_OUT, O 
                           => G_2665GAT_OUT);
   G_2664GAT : Nor_gate port map( I1 => G_2615GAT_OUT, I2 => G_2503GAT_OUT, O 
                           => G_2664GAT_OUT);
   G_2663GAT : Nor_gate port map( I1 => G_2564GAT_OUT, I2 => G_2615GAT_OUT, O 
                           => G_2663GAT_OUT);
   G_2662GAT : Nor_gate port map( I1 => G_2611GAT_OUT, I2 => G_2498GAT_OUT, O 
                           => G_2662GAT_OUT);
   G_2661GAT : Nor_gate port map( I1 => G_2561GAT_OUT, I2 => G_2611GAT_OUT, O 
                           => G_2661GAT_OUT);
   G_2660GAT : Nor_gate port map( I1 => G_2607GAT_OUT, I2 => G_2493GAT_OUT, O 
                           => G_2660GAT_OUT);
   G_2659GAT : Nor_gate port map( I1 => G_2558GAT_OUT, I2 => G_2607GAT_OUT, O 
                           => G_2659GAT_OUT);
   G_2658GAT : Nor_gate port map( I1 => G_2603GAT_OUT, I2 => G_2488GAT_OUT, O 
                           => G_2658GAT_OUT);
   G_2657GAT : Nor_gate port map( I1 => G_2555GAT_OUT, I2 => G_2603GAT_OUT, O 
                           => G_2657GAT_OUT);
   G_2656GAT : Nor_gate port map( I1 => G_2599GAT_OUT, I2 => G_2483GAT_OUT, O 
                           => G_2656GAT_OUT);
   G_2655GAT : Nor_gate port map( I1 => G_2552GAT_OUT, I2 => G_2599GAT_OUT, O 
                           => G_2655GAT_OUT);
   G_2654GAT : Nor_gate port map( I1 => G_2595GAT_OUT, I2 => G_2478GAT_OUT, O 
                           => G_2654GAT_OUT);
   G_2653GAT : Nor_gate port map( I1 => G_2549GAT_OUT, I2 => G_2595GAT_OUT, O 
                           => G_2653GAT_OUT);
   G_2650GAT : Nor_gate port map( I1 => G_2410GAT_OUT, I2 => G_2591GAT_OUT, O 
                           => G_2650GAT_OUT);
   G_2649GAT : Nor_gate port map( I1 => G_2591GAT_OUT, I2 => G_1230GAT_OUT, O 
                           => G_2649GAT_OUT);
   G_2648GAT : Nor_gate port map( I1 => G_2545GAT_OUT, I2 => G_2591GAT_OUT, O 
                           => G_2648GAT_OUT);
   G_2644GAT : Nor_gate port map( I1 => G_2588GAT_OUT, I2 => G_1182GAT_OUT, O 
                           => G_2644GAT_OUT);
   G_2641GAT : Nor_gate port map( I1 => G_2586GAT_OUT, I2 => G_2587GAT_OUT, O 
                           => G_2641GAT_OUT);
   G_2640GAT : Nor_gate port map( I1 => G_2582GAT_OUT, I2 => G_2533GAT_OUT, O 
                           => G_2640GAT_OUT);
   G_2639GAT : Nor_gate port map( I1 => G_2536GAT_OUT, I2 => G_2582GAT_OUT, O 
                           => G_2639GAT_OUT);
   G_2635GAT : Nor_gate port map( I1 => G_2579GAT_OUT, I2 => G_2528GAT_OUT, O 
                           => G_2635GAT_OUT);
   G_2631GAT : Nor_gate port map( I1 => G_2576GAT_OUT, I2 => G_2523GAT_OUT, O 
                           => G_2631GAT_OUT);
   G_2627GAT : Nor_gate port map( I1 => G_2573GAT_OUT, I2 => G_2518GAT_OUT, O 
                           => G_2627GAT_OUT);
   G_2623GAT : Nor_gate port map( I1 => G_2570GAT_OUT, I2 => G_2513GAT_OUT, O 
                           => G_2623GAT_OUT);
   G_2619GAT : Nor_gate port map( I1 => G_2567GAT_OUT, I2 => G_2508GAT_OUT, O 
                           => G_2619GAT_OUT);
   G_2615GAT : Nor_gate port map( I1 => G_2564GAT_OUT, I2 => G_2503GAT_OUT, O 
                           => G_2615GAT_OUT);
   G_2611GAT : Nor_gate port map( I1 => G_2561GAT_OUT, I2 => G_2498GAT_OUT, O 
                           => G_2611GAT_OUT);
   G_2607GAT : Nor_gate port map( I1 => G_2558GAT_OUT, I2 => G_2493GAT_OUT, O 
                           => G_2607GAT_OUT);
   G_2603GAT : Nor_gate port map( I1 => G_2555GAT_OUT, I2 => G_2488GAT_OUT, O 
                           => G_2603GAT_OUT);
   G_2599GAT : Nor_gate port map( I1 => G_2552GAT_OUT, I2 => G_2483GAT_OUT, O 
                           => G_2599GAT_OUT);
   G_2595GAT : Nor_gate port map( I1 => G_2549GAT_OUT, I2 => G_2478GAT_OUT, O 
                           => G_2595GAT_OUT);
   G_2591GAT : Nor_gate port map( I1 => G_2545GAT_OUT, I2 => G_1230GAT_OUT, O 
                           => G_2591GAT_OUT);
   G_2588GAT : Nor_gate port map( I1 => G_2543GAT_OUT, I2 => G_2544GAT_OUT, O 
                           => G_2588GAT_OUT);
   G_2587GAT : Nor_gate port map( I1 => G_2539GAT_OUT, I2 => G_2464GAT_OUT, O 
                           => G_2587GAT_OUT);
   G_2586GAT : Nor_gate port map( I1 => G_2467GAT_OUT, I2 => G_2539GAT_OUT, O 
                           => G_2586GAT_OUT);
   G_2582GAT : Nor_gate port map( I1 => G_2536GAT_OUT, I2 => G_2533GAT_OUT, O 
                           => G_2582GAT_OUT);
   G_2579GAT : Nor_gate port map( I1 => G_2531GAT_OUT, I2 => G_2532GAT_OUT, O 
                           => G_2579GAT_OUT);
   G_2576GAT : Nor_gate port map( I1 => G_2526GAT_OUT, I2 => G_2527GAT_OUT, O 
                           => G_2576GAT_OUT);
   G_2573GAT : Nor_gate port map( I1 => G_2521GAT_OUT, I2 => G_2522GAT_OUT, O 
                           => G_2573GAT_OUT);
   G_2570GAT : Nor_gate port map( I1 => G_2516GAT_OUT, I2 => G_2517GAT_OUT, O 
                           => G_2570GAT_OUT);
   G_2567GAT : Nor_gate port map( I1 => G_2511GAT_OUT, I2 => G_2512GAT_OUT, O 
                           => G_2567GAT_OUT);
   G_2564GAT : Nor_gate port map( I1 => G_2506GAT_OUT, I2 => G_2507GAT_OUT, O 
                           => G_2564GAT_OUT);
   G_2561GAT : Nor_gate port map( I1 => G_2501GAT_OUT, I2 => G_2502GAT_OUT, O 
                           => G_2561GAT_OUT);
   G_2558GAT : Nor_gate port map( I1 => G_2496GAT_OUT, I2 => G_2497GAT_OUT, O 
                           => G_2558GAT_OUT);
   G_2555GAT : Nor_gate port map( I1 => G_2491GAT_OUT, I2 => G_2492GAT_OUT, O 
                           => G_2555GAT_OUT);
   G_2552GAT : Nor_gate port map( I1 => G_2486GAT_OUT, I2 => G_2487GAT_OUT, O 
                           => G_2552GAT_OUT);
   G_2549GAT : Nor_gate port map( I1 => G_2481GAT_OUT, I2 => G_2482GAT_OUT, O 
                           => G_2549GAT_OUT);
   G_2545GAT : Nor_gate port map( I1 => G_2474GAT_OUT, I2 => G_2475GAT_OUT, O 
                           => G_2545GAT_OUT);
   G_2544GAT : Nor_gate port map( I1 => G_2470GAT_OUT, I2 => G_2404GAT_OUT, O 
                           => G_2544GAT_OUT);
   G_2543GAT : Nor_gate port map( I1 => G_2407GAT_OUT, I2 => G_2470GAT_OUT, O 
                           => G_2543GAT_OUT);
   G_2539GAT : Nor_gate port map( I1 => G_2467GAT_OUT, I2 => G_2464GAT_OUT, O 
                           => G_2539GAT_OUT);
   G_2536GAT : Nor_gate port map( I1 => G_2462GAT_OUT, I2 => G_2463GAT_OUT, O 
                           => G_2536GAT_OUT);
   G_2533GAT : Nor_gate port map( I1 => G_2313GAT_OUT, I2 => G_2458GAT_OUT, O 
                           => G_2533GAT_OUT);
   G_2532GAT : Nor_gate port map( I1 => G_2458GAT_OUT, I2 => G_1083GAT_OUT, O 
                           => G_2532GAT_OUT);
   G_2531GAT : Nor_gate port map( I1 => G_2395GAT_OUT, I2 => G_2458GAT_OUT, O 
                           => G_2531GAT_OUT);
   G_2528GAT : Nor_gate port map( I1 => G_2309GAT_OUT, I2 => G_2454GAT_OUT, O 
                           => G_2528GAT_OUT);
   G_2527GAT : Nor_gate port map( I1 => G_2454GAT_OUT, I2 => G_1035GAT_OUT, O 
                           => G_2527GAT_OUT);
   G_2526GAT : Nor_gate port map( I1 => G_2392GAT_OUT, I2 => G_2454GAT_OUT, O 
                           => G_2526GAT_OUT);
   G_2523GAT : Nor_gate port map( I1 => G_2305GAT_OUT, I2 => G_2450GAT_OUT, O 
                           => G_2523GAT_OUT);
   G_2522GAT : Nor_gate port map( I1 => G_2450GAT_OUT, I2 => G_987GAT_OUT, O =>
                           G_2522GAT_OUT);
   G_2521GAT : Nor_gate port map( I1 => G_2389GAT_OUT, I2 => G_2450GAT_OUT, O 
                           => G_2521GAT_OUT);
   G_2518GAT : Nor_gate port map( I1 => G_2301GAT_OUT, I2 => G_2446GAT_OUT, O 
                           => G_2518GAT_OUT);
   G_2517GAT : Nor_gate port map( I1 => G_2446GAT_OUT, I2 => G_939GAT_OUT, O =>
                           G_2517GAT_OUT);
   G_2516GAT : Nor_gate port map( I1 => G_2386GAT_OUT, I2 => G_2446GAT_OUT, O 
                           => G_2516GAT_OUT);
   G_2513GAT : Nor_gate port map( I1 => G_2297GAT_OUT, I2 => G_2442GAT_OUT, O 
                           => G_2513GAT_OUT);
   G_2512GAT : Nor_gate port map( I1 => G_2442GAT_OUT, I2 => G_891GAT_OUT, O =>
                           G_2512GAT_OUT);
   G_2511GAT : Nor_gate port map( I1 => G_2383GAT_OUT, I2 => G_2442GAT_OUT, O 
                           => G_2511GAT_OUT);
   G_2508GAT : Nor_gate port map( I1 => G_2293GAT_OUT, I2 => G_2438GAT_OUT, O 
                           => G_2508GAT_OUT);
   G_2507GAT : Nor_gate port map( I1 => G_2438GAT_OUT, I2 => G_843GAT_OUT, O =>
                           G_2507GAT_OUT);
   G_2506GAT : Nor_gate port map( I1 => G_2380GAT_OUT, I2 => G_2438GAT_OUT, O 
                           => G_2506GAT_OUT);
   G_2503GAT : Nor_gate port map( I1 => G_2289GAT_OUT, I2 => G_2434GAT_OUT, O 
                           => G_2503GAT_OUT);
   G_2502GAT : Nor_gate port map( I1 => G_2434GAT_OUT, I2 => G_795GAT_OUT, O =>
                           G_2502GAT_OUT);
   G_2501GAT : Nor_gate port map( I1 => G_2377GAT_OUT, I2 => G_2434GAT_OUT, O 
                           => G_2501GAT_OUT);
   G_2498GAT : Nor_gate port map( I1 => G_2285GAT_OUT, I2 => G_2430GAT_OUT, O 
                           => G_2498GAT_OUT);
   G_2497GAT : Nor_gate port map( I1 => G_2430GAT_OUT, I2 => G_747GAT_OUT, O =>
                           G_2497GAT_OUT);
   G_2496GAT : Nor_gate port map( I1 => G_2374GAT_OUT, I2 => G_2430GAT_OUT, O 
                           => G_2496GAT_OUT);
   G_2493GAT : Nor_gate port map( I1 => G_2281GAT_OUT, I2 => G_2426GAT_OUT, O 
                           => G_2493GAT_OUT);
   G_2492GAT : Nor_gate port map( I1 => G_2426GAT_OUT, I2 => G_699GAT_OUT, O =>
                           G_2492GAT_OUT);
   G_2491GAT : Nor_gate port map( I1 => G_2371GAT_OUT, I2 => G_2426GAT_OUT, O 
                           => G_2491GAT_OUT);
   G_2488GAT : Nor_gate port map( I1 => G_2277GAT_OUT, I2 => G_2422GAT_OUT, O 
                           => G_2488GAT_OUT);
   G_2487GAT : Nor_gate port map( I1 => G_2422GAT_OUT, I2 => G_651GAT_OUT, O =>
                           G_2487GAT_OUT);
   G_2486GAT : Nor_gate port map( I1 => G_2368GAT_OUT, I2 => G_2422GAT_OUT, O 
                           => G_2486GAT_OUT);
   G_2483GAT : Nor_gate port map( I1 => G_2273GAT_OUT, I2 => G_2418GAT_OUT, O 
                           => G_2483GAT_OUT);
   G_2482GAT : Nor_gate port map( I1 => G_2418GAT_OUT, I2 => G_603GAT_OUT, O =>
                           G_2482GAT_OUT);
   G_2481GAT : Nor_gate port map( I1 => G_2365GAT_OUT, I2 => G_2418GAT_OUT, O 
                           => G_2481GAT_OUT);
   G_2478GAT : Nor_gate port map( I1 => G_2269GAT_OUT, I2 => G_2414GAT_OUT, O 
                           => G_2478GAT_OUT);
   G_2477GAT : Nor_gate port map( I1 => G_2414GAT_OUT, I2 => G_555GAT_OUT, O =>
                           G_2477GAT_OUT);
   G_2476GAT : Nor_gate port map( I1 => G_2362GAT_OUT, I2 => G_2414GAT_OUT, O 
                           => G_2476GAT_OUT);
   G_2475GAT : Nor_gate port map( I1 => G_2410GAT_OUT, I2 => G_2359GAT_OUT, O 
                           => G_2475GAT_OUT);
   G_2474GAT : Nor_gate port map( I1 => G_1275GAT_OUT, I2 => G_2410GAT_OUT, O 
                           => G_2474GAT_OUT);
   G_2470GAT : Nor_gate port map( I1 => G_2407GAT_OUT, I2 => G_2404GAT_OUT, O 
                           => G_2470GAT_OUT);
   G_2467GAT : Nor_gate port map( I1 => G_2402GAT_OUT, I2 => G_2403GAT_OUT, O 
                           => G_2467GAT_OUT);
   G_2464GAT : Nor_gate port map( I1 => G_2260GAT_OUT, I2 => G_2398GAT_OUT, O 
                           => G_2464GAT_OUT);
   G_2463GAT : Nor_gate port map( I1 => G_2398GAT_OUT, I2 => G_1131GAT_OUT, O 
                           => G_2463GAT_OUT);
   G_2462GAT : Nor_gate port map( I1 => G_2350GAT_OUT, I2 => G_2398GAT_OUT, O 
                           => G_2462GAT_OUT);
   G_2458GAT : Nor_gate port map( I1 => G_2395GAT_OUT, I2 => G_1083GAT_OUT, O 
                           => G_2458GAT_OUT);
   G_2454GAT : Nor_gate port map( I1 => G_2392GAT_OUT, I2 => G_1035GAT_OUT, O 
                           => G_2454GAT_OUT);
   G_2450GAT : Nor_gate port map( I1 => G_2389GAT_OUT, I2 => G_987GAT_OUT, O =>
                           G_2450GAT_OUT);
   G_2446GAT : Nor_gate port map( I1 => G_2386GAT_OUT, I2 => G_939GAT_OUT, O =>
                           G_2446GAT_OUT);
   G_2442GAT : Nor_gate port map( I1 => G_2383GAT_OUT, I2 => G_891GAT_OUT, O =>
                           G_2442GAT_OUT);
   G_2438GAT : Nor_gate port map( I1 => G_2380GAT_OUT, I2 => G_843GAT_OUT, O =>
                           G_2438GAT_OUT);
   G_2434GAT : Nor_gate port map( I1 => G_2377GAT_OUT, I2 => G_795GAT_OUT, O =>
                           G_2434GAT_OUT);
   G_2430GAT : Nor_gate port map( I1 => G_2374GAT_OUT, I2 => G_747GAT_OUT, O =>
                           G_2430GAT_OUT);
   G_2426GAT : Nor_gate port map( I1 => G_2371GAT_OUT, I2 => G_699GAT_OUT, O =>
                           G_2426GAT_OUT);
   G_2422GAT : Nor_gate port map( I1 => G_2368GAT_OUT, I2 => G_651GAT_OUT, O =>
                           G_2422GAT_OUT);
   G_2418GAT : Nor_gate port map( I1 => G_2365GAT_OUT, I2 => G_603GAT_OUT, O =>
                           G_2418GAT_OUT);
   G_2414GAT : Nor_gate port map( I1 => G_2362GAT_OUT, I2 => G_555GAT_OUT, O =>
                           G_2414GAT_OUT);
   G_2410GAT : Nor_gate port map( I1 => G_1275GAT_OUT, I2 => G_2359GAT_OUT, O 
                           => G_2410GAT_OUT);
   G_2407GAT : Nor_gate port map( I1 => G_2357GAT_OUT, I2 => G_2358GAT_OUT, O 
                           => G_2407GAT_OUT);
   G_2404GAT : Nor_gate port map( I1 => G_2217GAT_OUT, I2 => G_2353GAT_OUT, O 
                           => G_2404GAT_OUT);
   G_2403GAT : Nor_gate port map( I1 => G_2353GAT_OUT, I2 => G_1179GAT_OUT, O 
                           => G_2403GAT_OUT);
   G_2402GAT : Nor_gate port map( I1 => G_2319GAT_OUT, I2 => G_2353GAT_OUT, O 
                           => G_2402GAT_OUT);
   G_2398GAT : Nor_gate port map( I1 => G_2350GAT_OUT, I2 => G_1131GAT_OUT, O 
                           => G_2398GAT_OUT);
   G_2395GAT : Nor_gate port map( I1 => G_2348GAT_OUT, I2 => G_2349GAT_OUT, O 
                           => G_2395GAT_OUT);
   G_2392GAT : Nor_gate port map( I1 => G_2346GAT_OUT, I2 => G_2347GAT_OUT, O 
                           => G_2392GAT_OUT);
   G_2389GAT : Nor_gate port map( I1 => G_2344GAT_OUT, I2 => G_2345GAT_OUT, O 
                           => G_2389GAT_OUT);
   G_2386GAT : Nor_gate port map( I1 => G_2342GAT_OUT, I2 => G_2343GAT_OUT, O 
                           => G_2386GAT_OUT);
   G_2383GAT : Nor_gate port map( I1 => G_2340GAT_OUT, I2 => G_2341GAT_OUT, O 
                           => G_2383GAT_OUT);
   G_2380GAT : Nor_gate port map( I1 => G_2338GAT_OUT, I2 => G_2339GAT_OUT, O 
                           => G_2380GAT_OUT);
   G_2377GAT : Nor_gate port map( I1 => G_2336GAT_OUT, I2 => G_2337GAT_OUT, O 
                           => G_2377GAT_OUT);
   G_2374GAT : Nor_gate port map( I1 => G_2334GAT_OUT, I2 => G_2335GAT_OUT, O 
                           => G_2374GAT_OUT);
   G_2371GAT : Nor_gate port map( I1 => G_2332GAT_OUT, I2 => G_2333GAT_OUT, O 
                           => G_2371GAT_OUT);
   G_2368GAT : Nor_gate port map( I1 => G_2330GAT_OUT, I2 => G_2331GAT_OUT, O 
                           => G_2368GAT_OUT);
   G_2365GAT : Nor_gate port map( I1 => G_2328GAT_OUT, I2 => G_2329GAT_OUT, O 
                           => G_2365GAT_OUT);
   G_2362GAT : Nor_gate port map( I1 => G_2326GAT_OUT, I2 => G_2327GAT_OUT, O 
                           => G_2362GAT_OUT);
   G_2359GAT : Nor_gate port map( I1 => G_2145GAT_OUT, I2 => G_2322GAT_OUT, O 
                           => G_2359GAT_OUT);
   G_2358GAT : Nor_gate port map( I1 => G_2322GAT_OUT, I2 => G_1227GAT_OUT, O 
                           => G_2358GAT_OUT);
   G_2357GAT : Nor_gate port map( I1 => G_2266GAT_OUT, I2 => G_2322GAT_OUT, O 
                           => G_2357GAT_OUT);
   G_2353GAT : Nor_gate port map( I1 => G_2319GAT_OUT, I2 => G_1179GAT_OUT, O 
                           => G_2353GAT_OUT);
   G_2350GAT : Nor_gate port map( I1 => G_2317GAT_OUT, I2 => G_2318GAT_OUT, O 
                           => G_2350GAT_OUT);
   G_2349GAT : Nor_gate port map( I1 => G_2313GAT_OUT, I2 => G_2206GAT_OUT, O 
                           => G_2349GAT_OUT);
   G_2348GAT : Nor_gate port map( I1 => G_2257GAT_OUT, I2 => G_2313GAT_OUT, O 
                           => G_2348GAT_OUT);
   G_2347GAT : Nor_gate port map( I1 => G_2309GAT_OUT, I2 => G_2201GAT_OUT, O 
                           => G_2347GAT_OUT);
   G_2346GAT : Nor_gate port map( I1 => G_2254GAT_OUT, I2 => G_2309GAT_OUT, O 
                           => G_2346GAT_OUT);
   G_2345GAT : Nor_gate port map( I1 => G_2305GAT_OUT, I2 => G_2196GAT_OUT, O 
                           => G_2345GAT_OUT);
   G_2344GAT : Nor_gate port map( I1 => G_2251GAT_OUT, I2 => G_2305GAT_OUT, O 
                           => G_2344GAT_OUT);
   G_2343GAT : Nor_gate port map( I1 => G_2301GAT_OUT, I2 => G_2191GAT_OUT, O 
                           => G_2343GAT_OUT);
   G_2342GAT : Nor_gate port map( I1 => G_2248GAT_OUT, I2 => G_2301GAT_OUT, O 
                           => G_2342GAT_OUT);
   G_2341GAT : Nor_gate port map( I1 => G_2297GAT_OUT, I2 => G_2186GAT_OUT, O 
                           => G_2341GAT_OUT);
   G_2340GAT : Nor_gate port map( I1 => G_2245GAT_OUT, I2 => G_2297GAT_OUT, O 
                           => G_2340GAT_OUT);
   G_2339GAT : Nor_gate port map( I1 => G_2293GAT_OUT, I2 => G_2181GAT_OUT, O 
                           => G_2339GAT_OUT);
   G_2338GAT : Nor_gate port map( I1 => G_2242GAT_OUT, I2 => G_2293GAT_OUT, O 
                           => G_2338GAT_OUT);
   G_2337GAT : Nor_gate port map( I1 => G_2289GAT_OUT, I2 => G_2176GAT_OUT, O 
                           => G_2337GAT_OUT);
   G_2336GAT : Nor_gate port map( I1 => G_2239GAT_OUT, I2 => G_2289GAT_OUT, O 
                           => G_2336GAT_OUT);
   G_2335GAT : Nor_gate port map( I1 => G_2285GAT_OUT, I2 => G_2171GAT_OUT, O 
                           => G_2335GAT_OUT);
   G_2334GAT : Nor_gate port map( I1 => G_2236GAT_OUT, I2 => G_2285GAT_OUT, O 
                           => G_2334GAT_OUT);
   G_2333GAT : Nor_gate port map( I1 => G_2281GAT_OUT, I2 => G_2166GAT_OUT, O 
                           => G_2333GAT_OUT);
   G_2332GAT : Nor_gate port map( I1 => G_2233GAT_OUT, I2 => G_2281GAT_OUT, O 
                           => G_2332GAT_OUT);
   G_2331GAT : Nor_gate port map( I1 => G_2277GAT_OUT, I2 => G_2161GAT_OUT, O 
                           => G_2331GAT_OUT);
   G_2330GAT : Nor_gate port map( I1 => G_2230GAT_OUT, I2 => G_2277GAT_OUT, O 
                           => G_2330GAT_OUT);
   G_2329GAT : Nor_gate port map( I1 => G_2273GAT_OUT, I2 => G_2156GAT_OUT, O 
                           => G_2329GAT_OUT);
   G_2328GAT : Nor_gate port map( I1 => G_2227GAT_OUT, I2 => G_2273GAT_OUT, O 
                           => G_2328GAT_OUT);
   G_2327GAT : Nor_gate port map( I1 => G_2269GAT_OUT, I2 => G_2151GAT_OUT, O 
                           => G_2327GAT_OUT);
   G_2326GAT : Nor_gate port map( I1 => G_2224GAT_OUT, I2 => G_2269GAT_OUT, O 
                           => G_2326GAT_OUT);
   G_2322GAT : Nor_gate port map( I1 => G_2266GAT_OUT, I2 => G_1227GAT_OUT, O 
                           => G_2322GAT_OUT);
   G_2319GAT : Nor_gate port map( I1 => G_2264GAT_OUT, I2 => G_2265GAT_OUT, O 
                           => G_2319GAT_OUT);
   G_2318GAT : Nor_gate port map( I1 => G_2260GAT_OUT, I2 => G_2211GAT_OUT, O 
                           => G_2318GAT_OUT);
   G_2317GAT : Nor_gate port map( I1 => G_2214GAT_OUT, I2 => G_2260GAT_OUT, O 
                           => G_2317GAT_OUT);
   G_2313GAT : Nor_gate port map( I1 => G_2257GAT_OUT, I2 => G_2206GAT_OUT, O 
                           => G_2313GAT_OUT);
   G_2309GAT : Nor_gate port map( I1 => G_2254GAT_OUT, I2 => G_2201GAT_OUT, O 
                           => G_2309GAT_OUT);
   G_2305GAT : Nor_gate port map( I1 => G_2251GAT_OUT, I2 => G_2196GAT_OUT, O 
                           => G_2305GAT_OUT);
   G_2301GAT : Nor_gate port map( I1 => G_2248GAT_OUT, I2 => G_2191GAT_OUT, O 
                           => G_2301GAT_OUT);
   G_2297GAT : Nor_gate port map( I1 => G_2245GAT_OUT, I2 => G_2186GAT_OUT, O 
                           => G_2297GAT_OUT);
   G_2293GAT : Nor_gate port map( I1 => G_2242GAT_OUT, I2 => G_2181GAT_OUT, O 
                           => G_2293GAT_OUT);
   G_2289GAT : Nor_gate port map( I1 => G_2239GAT_OUT, I2 => G_2176GAT_OUT, O 
                           => G_2289GAT_OUT);
   G_2285GAT : Nor_gate port map( I1 => G_2236GAT_OUT, I2 => G_2171GAT_OUT, O 
                           => G_2285GAT_OUT);
   G_2281GAT : Nor_gate port map( I1 => G_2233GAT_OUT, I2 => G_2166GAT_OUT, O 
                           => G_2281GAT_OUT);
   G_2277GAT : Nor_gate port map( I1 => G_2230GAT_OUT, I2 => G_2161GAT_OUT, O 
                           => G_2277GAT_OUT);
   G_2273GAT : Nor_gate port map( I1 => G_2227GAT_OUT, I2 => G_2156GAT_OUT, O 
                           => G_2273GAT_OUT);
   G_2269GAT : Nor_gate port map( I1 => G_2224GAT_OUT, I2 => G_2151GAT_OUT, O 
                           => G_2269GAT_OUT);
   G_2266GAT : Nor_gate port map( I1 => G_2221GAT_OUT, I2 => G_2222GAT_OUT, O 
                           => G_2266GAT_OUT);
   G_2265GAT : Nor_gate port map( I1 => G_2217GAT_OUT, I2 => G_2139GAT_OUT, O 
                           => G_2265GAT_OUT);
   G_2264GAT : Nor_gate port map( I1 => G_2142GAT_OUT, I2 => G_2217GAT_OUT, O 
                           => G_2264GAT_OUT);
   G_2260GAT : Nor_gate port map( I1 => G_2214GAT_OUT, I2 => G_2211GAT_OUT, O 
                           => G_2260GAT_OUT);
   G_2257GAT : Nor_gate port map( I1 => G_2209GAT_OUT, I2 => G_2210GAT_OUT, O 
                           => G_2257GAT_OUT);
   G_2254GAT : Nor_gate port map( I1 => G_2204GAT_OUT, I2 => G_2205GAT_OUT, O 
                           => G_2254GAT_OUT);
   G_2251GAT : Nor_gate port map( I1 => G_2199GAT_OUT, I2 => G_2200GAT_OUT, O 
                           => G_2251GAT_OUT);
   G_2248GAT : Nor_gate port map( I1 => G_2194GAT_OUT, I2 => G_2195GAT_OUT, O 
                           => G_2248GAT_OUT);
   G_2245GAT : Nor_gate port map( I1 => G_2189GAT_OUT, I2 => G_2190GAT_OUT, O 
                           => G_2245GAT_OUT);
   G_2242GAT : Nor_gate port map( I1 => G_2184GAT_OUT, I2 => G_2185GAT_OUT, O 
                           => G_2242GAT_OUT);
   G_2239GAT : Nor_gate port map( I1 => G_2179GAT_OUT, I2 => G_2180GAT_OUT, O 
                           => G_2239GAT_OUT);
   G_2236GAT : Nor_gate port map( I1 => G_2174GAT_OUT, I2 => G_2175GAT_OUT, O 
                           => G_2236GAT_OUT);
   G_2233GAT : Nor_gate port map( I1 => G_2169GAT_OUT, I2 => G_2170GAT_OUT, O 
                           => G_2233GAT_OUT);
   G_2230GAT : Nor_gate port map( I1 => G_2164GAT_OUT, I2 => G_2165GAT_OUT, O 
                           => G_2230GAT_OUT);
   G_2227GAT : Nor_gate port map( I1 => G_2159GAT_OUT, I2 => G_2160GAT_OUT, O 
                           => G_2227GAT_OUT);
   G_2224GAT : Nor_gate port map( I1 => G_2154GAT_OUT, I2 => G_2155GAT_OUT, O 
                           => G_2224GAT_OUT);
   G_2222GAT : Nor_gate port map( I1 => G_2145GAT_OUT, I2 => G_2082GAT_OUT, O 
                           => G_2222GAT_OUT);
   G_2221GAT : Nor_gate port map( I1 => G_1272GAT_OUT, I2 => G_2145GAT_OUT, O 
                           => G_2221GAT_OUT);
   G_2217GAT : Nor_gate port map( I1 => G_2142GAT_OUT, I2 => G_2139GAT_OUT, O 
                           => G_2217GAT_OUT);
   G_2214GAT : Nor_gate port map( I1 => G_2137GAT_OUT, I2 => G_2138GAT_OUT, O 
                           => G_2214GAT_OUT);
   G_2211GAT : Nor_gate port map( I1 => G_1995GAT_OUT, I2 => G_2133GAT_OUT, O 
                           => G_2211GAT_OUT);
   G_2210GAT : Nor_gate port map( I1 => G_2133GAT_OUT, I2 => G_1128GAT_OUT, O 
                           => G_2210GAT_OUT);
   G_2209GAT : Nor_gate port map( I1 => G_2073GAT_OUT, I2 => G_2133GAT_OUT, O 
                           => G_2209GAT_OUT);
   G_2206GAT : Nor_gate port map( I1 => G_1991GAT_OUT, I2 => G_2129GAT_OUT, O 
                           => G_2206GAT_OUT);
   G_2205GAT : Nor_gate port map( I1 => G_2129GAT_OUT, I2 => G_1080GAT_OUT, O 
                           => G_2205GAT_OUT);
   G_2204GAT : Nor_gate port map( I1 => G_2070GAT_OUT, I2 => G_2129GAT_OUT, O 
                           => G_2204GAT_OUT);
   G_2201GAT : Nor_gate port map( I1 => G_1987GAT_OUT, I2 => G_2125GAT_OUT, O 
                           => G_2201GAT_OUT);
   G_2200GAT : Nor_gate port map( I1 => G_2125GAT_OUT, I2 => G_1032GAT_OUT, O 
                           => G_2200GAT_OUT);
   G_2199GAT : Nor_gate port map( I1 => G_2067GAT_OUT, I2 => G_2125GAT_OUT, O 
                           => G_2199GAT_OUT);
   G_2196GAT : Nor_gate port map( I1 => G_1983GAT_OUT, I2 => G_2121GAT_OUT, O 
                           => G_2196GAT_OUT);
   G_2195GAT : Nor_gate port map( I1 => G_2121GAT_OUT, I2 => G_984GAT_OUT, O =>
                           G_2195GAT_OUT);
   G_2194GAT : Nor_gate port map( I1 => G_2064GAT_OUT, I2 => G_2121GAT_OUT, O 
                           => G_2194GAT_OUT);
   G_2191GAT : Nor_gate port map( I1 => G_1979GAT_OUT, I2 => G_2117GAT_OUT, O 
                           => G_2191GAT_OUT);
   G_2190GAT : Nor_gate port map( I1 => G_2117GAT_OUT, I2 => G_936GAT_OUT, O =>
                           G_2190GAT_OUT);
   G_2189GAT : Nor_gate port map( I1 => G_2061GAT_OUT, I2 => G_2117GAT_OUT, O 
                           => G_2189GAT_OUT);
   G_2186GAT : Nor_gate port map( I1 => G_1975GAT_OUT, I2 => G_2113GAT_OUT, O 
                           => G_2186GAT_OUT);
   G_2185GAT : Nor_gate port map( I1 => G_2113GAT_OUT, I2 => G_888GAT_OUT, O =>
                           G_2185GAT_OUT);
   G_2184GAT : Nor_gate port map( I1 => G_2058GAT_OUT, I2 => G_2113GAT_OUT, O 
                           => G_2184GAT_OUT);
   G_2181GAT : Nor_gate port map( I1 => G_1971GAT_OUT, I2 => G_2109GAT_OUT, O 
                           => G_2181GAT_OUT);
   G_2180GAT : Nor_gate port map( I1 => G_2109GAT_OUT, I2 => G_840GAT_OUT, O =>
                           G_2180GAT_OUT);
   G_2179GAT : Nor_gate port map( I1 => G_2055GAT_OUT, I2 => G_2109GAT_OUT, O 
                           => G_2179GAT_OUT);
   G_2176GAT : Nor_gate port map( I1 => G_1967GAT_OUT, I2 => G_2105GAT_OUT, O 
                           => G_2176GAT_OUT);
   G_2175GAT : Nor_gate port map( I1 => G_2105GAT_OUT, I2 => G_792GAT_OUT, O =>
                           G_2175GAT_OUT);
   G_2174GAT : Nor_gate port map( I1 => G_2052GAT_OUT, I2 => G_2105GAT_OUT, O 
                           => G_2174GAT_OUT);
   G_2171GAT : Nor_gate port map( I1 => G_1963GAT_OUT, I2 => G_2101GAT_OUT, O 
                           => G_2171GAT_OUT);
   G_2170GAT : Nor_gate port map( I1 => G_2101GAT_OUT, I2 => G_744GAT_OUT, O =>
                           G_2170GAT_OUT);
   G_2169GAT : Nor_gate port map( I1 => G_2049GAT_OUT, I2 => G_2101GAT_OUT, O 
                           => G_2169GAT_OUT);
   G_2166GAT : Nor_gate port map( I1 => G_1959GAT_OUT, I2 => G_2097GAT_OUT, O 
                           => G_2166GAT_OUT);
   G_2165GAT : Nor_gate port map( I1 => G_2097GAT_OUT, I2 => G_696GAT_OUT, O =>
                           G_2165GAT_OUT);
   G_2164GAT : Nor_gate port map( I1 => G_2046GAT_OUT, I2 => G_2097GAT_OUT, O 
                           => G_2164GAT_OUT);
   G_2161GAT : Nor_gate port map( I1 => G_1955GAT_OUT, I2 => G_2093GAT_OUT, O 
                           => G_2161GAT_OUT);
   G_2160GAT : Nor_gate port map( I1 => G_2093GAT_OUT, I2 => G_648GAT_OUT, O =>
                           G_2160GAT_OUT);
   G_2159GAT : Nor_gate port map( I1 => G_2043GAT_OUT, I2 => G_2093GAT_OUT, O 
                           => G_2159GAT_OUT);
   G_2156GAT : Nor_gate port map( I1 => G_1951GAT_OUT, I2 => G_2089GAT_OUT, O 
                           => G_2156GAT_OUT);
   G_2155GAT : Nor_gate port map( I1 => G_2089GAT_OUT, I2 => G_600GAT_OUT, O =>
                           G_2155GAT_OUT);
   G_2154GAT : Nor_gate port map( I1 => G_2040GAT_OUT, I2 => G_2089GAT_OUT, O 
                           => G_2154GAT_OUT);
   G_2151GAT : Nor_gate port map( I1 => G_1947GAT_OUT, I2 => G_2085GAT_OUT, O 
                           => G_2151GAT_OUT);
   G_2150GAT : Nor_gate port map( I1 => G_2085GAT_OUT, I2 => G_552GAT_OUT, O =>
                           G_2150GAT_OUT);
   G_2149GAT : Nor_gate port map( I1 => G_2037GAT_OUT, I2 => G_2085GAT_OUT, O 
                           => G_2149GAT_OUT);
   G_2145GAT : Nor_gate port map( I1 => G_1272GAT_OUT, I2 => G_2082GAT_OUT, O 
                           => G_2145GAT_OUT);
   G_2142GAT : Nor_gate port map( I1 => G_2080GAT_OUT, I2 => G_2081GAT_OUT, O 
                           => G_2142GAT_OUT);
   G_2139GAT : Nor_gate port map( I1 => G_1941GAT_OUT, I2 => G_2076GAT_OUT, O 
                           => G_2139GAT_OUT);
   G_2138GAT : Nor_gate port map( I1 => G_2076GAT_OUT, I2 => G_1176GAT_OUT, O 
                           => G_2138GAT_OUT);
   G_2137GAT : Nor_gate port map( I1 => G_2030GAT_OUT, I2 => G_2076GAT_OUT, O 
                           => G_2137GAT_OUT);
   G_2133GAT : Nor_gate port map( I1 => G_2073GAT_OUT, I2 => G_1128GAT_OUT, O 
                           => G_2133GAT_OUT);
   G_2129GAT : Nor_gate port map( I1 => G_2070GAT_OUT, I2 => G_1080GAT_OUT, O 
                           => G_2129GAT_OUT);
   G_2125GAT : Nor_gate port map( I1 => G_2067GAT_OUT, I2 => G_1032GAT_OUT, O 
                           => G_2125GAT_OUT);
   G_2121GAT : Nor_gate port map( I1 => G_2064GAT_OUT, I2 => G_984GAT_OUT, O =>
                           G_2121GAT_OUT);
   G_2117GAT : Nor_gate port map( I1 => G_2061GAT_OUT, I2 => G_936GAT_OUT, O =>
                           G_2117GAT_OUT);
   G_2113GAT : Nor_gate port map( I1 => G_2058GAT_OUT, I2 => G_888GAT_OUT, O =>
                           G_2113GAT_OUT);
   G_2109GAT : Nor_gate port map( I1 => G_2055GAT_OUT, I2 => G_840GAT_OUT, O =>
                           G_2109GAT_OUT);
   G_2105GAT : Nor_gate port map( I1 => G_2052GAT_OUT, I2 => G_792GAT_OUT, O =>
                           G_2105GAT_OUT);
   G_2101GAT : Nor_gate port map( I1 => G_2049GAT_OUT, I2 => G_744GAT_OUT, O =>
                           G_2101GAT_OUT);
   G_2097GAT : Nor_gate port map( I1 => G_2046GAT_OUT, I2 => G_696GAT_OUT, O =>
                           G_2097GAT_OUT);
   G_2093GAT : Nor_gate port map( I1 => G_2043GAT_OUT, I2 => G_648GAT_OUT, O =>
                           G_2093GAT_OUT);
   G_2089GAT : Nor_gate port map( I1 => G_2040GAT_OUT, I2 => G_600GAT_OUT, O =>
                           G_2089GAT_OUT);
   G_2085GAT : Nor_gate port map( I1 => G_2037GAT_OUT, I2 => G_552GAT_OUT, O =>
                           G_2085GAT_OUT);
   G_2082GAT : Nor_gate port map( I1 => G_1897GAT_OUT, I2 => G_2033GAT_OUT, O 
                           => G_2082GAT_OUT);
   G_2081GAT : Nor_gate port map( I1 => G_2033GAT_OUT, I2 => G_1224GAT_OUT, O 
                           => G_2081GAT_OUT);
   G_2080GAT : Nor_gate port map( I1 => G_2001GAT_OUT, I2 => G_2033GAT_OUT, O 
                           => G_2080GAT_OUT);
   G_2076GAT : Nor_gate port map( I1 => G_2030GAT_OUT, I2 => G_1176GAT_OUT, O 
                           => G_2076GAT_OUT);
   G_2073GAT : Nor_gate port map( I1 => G_2028GAT_OUT, I2 => G_2029GAT_OUT, O 
                           => G_2073GAT_OUT);
   G_2070GAT : Nor_gate port map( I1 => G_2026GAT_OUT, I2 => G_2027GAT_OUT, O 
                           => G_2070GAT_OUT);
   G_2067GAT : Nor_gate port map( I1 => G_2024GAT_OUT, I2 => G_2025GAT_OUT, O 
                           => G_2067GAT_OUT);
   G_2064GAT : Nor_gate port map( I1 => G_2022GAT_OUT, I2 => G_2023GAT_OUT, O 
                           => G_2064GAT_OUT);
   G_2061GAT : Nor_gate port map( I1 => G_2020GAT_OUT, I2 => G_2021GAT_OUT, O 
                           => G_2061GAT_OUT);
   G_2058GAT : Nor_gate port map( I1 => G_2018GAT_OUT, I2 => G_2019GAT_OUT, O 
                           => G_2058GAT_OUT);
   G_2055GAT : Nor_gate port map( I1 => G_2016GAT_OUT, I2 => G_2017GAT_OUT, O 
                           => G_2055GAT_OUT);
   G_2052GAT : Nor_gate port map( I1 => G_2014GAT_OUT, I2 => G_2015GAT_OUT, O 
                           => G_2052GAT_OUT);
   G_2049GAT : Nor_gate port map( I1 => G_2012GAT_OUT, I2 => G_2013GAT_OUT, O 
                           => G_2049GAT_OUT);
   G_2046GAT : Nor_gate port map( I1 => G_2010GAT_OUT, I2 => G_2011GAT_OUT, O 
                           => G_2046GAT_OUT);
   G_2043GAT : Nor_gate port map( I1 => G_2008GAT_OUT, I2 => G_2009GAT_OUT, O 
                           => G_2043GAT_OUT);
   G_2040GAT : Nor_gate port map( I1 => G_2006GAT_OUT, I2 => G_2007GAT_OUT, O 
                           => G_2040GAT_OUT);
   G_2037GAT : Nor_gate port map( I1 => G_2004GAT_OUT, I2 => G_2005GAT_OUT, O 
                           => G_2037GAT_OUT);
   G_2033GAT : Nor_gate port map( I1 => G_2001GAT_OUT, I2 => G_1224GAT_OUT, O 
                           => G_2033GAT_OUT);
   G_2030GAT : Nor_gate port map( I1 => G_1999GAT_OUT, I2 => G_2000GAT_OUT, O 
                           => G_2030GAT_OUT);
   G_2029GAT : Nor_gate port map( I1 => G_1995GAT_OUT, I2 => G_1886GAT_OUT, O 
                           => G_2029GAT_OUT);
   G_2028GAT : Nor_gate port map( I1 => G_1938GAT_OUT, I2 => G_1995GAT_OUT, O 
                           => G_2028GAT_OUT);
   G_2027GAT : Nor_gate port map( I1 => G_1991GAT_OUT, I2 => G_1881GAT_OUT, O 
                           => G_2027GAT_OUT);
   G_2026GAT : Nor_gate port map( I1 => G_1935GAT_OUT, I2 => G_1991GAT_OUT, O 
                           => G_2026GAT_OUT);
   G_2025GAT : Nor_gate port map( I1 => G_1987GAT_OUT, I2 => G_1876GAT_OUT, O 
                           => G_2025GAT_OUT);
   G_2024GAT : Nor_gate port map( I1 => G_1932GAT_OUT, I2 => G_1987GAT_OUT, O 
                           => G_2024GAT_OUT);
   G_2023GAT : Nor_gate port map( I1 => G_1983GAT_OUT, I2 => G_1871GAT_OUT, O 
                           => G_2023GAT_OUT);
   G_2022GAT : Nor_gate port map( I1 => G_1929GAT_OUT, I2 => G_1983GAT_OUT, O 
                           => G_2022GAT_OUT);
   G_2021GAT : Nor_gate port map( I1 => G_1979GAT_OUT, I2 => G_1866GAT_OUT, O 
                           => G_2021GAT_OUT);
   G_2020GAT : Nor_gate port map( I1 => G_1926GAT_OUT, I2 => G_1979GAT_OUT, O 
                           => G_2020GAT_OUT);
   G_2019GAT : Nor_gate port map( I1 => G_1975GAT_OUT, I2 => G_1861GAT_OUT, O 
                           => G_2019GAT_OUT);
   G_2018GAT : Nor_gate port map( I1 => G_1923GAT_OUT, I2 => G_1975GAT_OUT, O 
                           => G_2018GAT_OUT);
   G_2017GAT : Nor_gate port map( I1 => G_1971GAT_OUT, I2 => G_1856GAT_OUT, O 
                           => G_2017GAT_OUT);
   G_2016GAT : Nor_gate port map( I1 => G_1920GAT_OUT, I2 => G_1971GAT_OUT, O 
                           => G_2016GAT_OUT);
   G_2015GAT : Nor_gate port map( I1 => G_1967GAT_OUT, I2 => G_1851GAT_OUT, O 
                           => G_2015GAT_OUT);
   G_2014GAT : Nor_gate port map( I1 => G_1917GAT_OUT, I2 => G_1967GAT_OUT, O 
                           => G_2014GAT_OUT);
   G_2013GAT : Nor_gate port map( I1 => G_1963GAT_OUT, I2 => G_1846GAT_OUT, O 
                           => G_2013GAT_OUT);
   G_2012GAT : Nor_gate port map( I1 => G_1914GAT_OUT, I2 => G_1963GAT_OUT, O 
                           => G_2012GAT_OUT);
   G_2011GAT : Nor_gate port map( I1 => G_1959GAT_OUT, I2 => G_1841GAT_OUT, O 
                           => G_2011GAT_OUT);
   G_2010GAT : Nor_gate port map( I1 => G_1911GAT_OUT, I2 => G_1959GAT_OUT, O 
                           => G_2010GAT_OUT);
   G_2009GAT : Nor_gate port map( I1 => G_1955GAT_OUT, I2 => G_1836GAT_OUT, O 
                           => G_2009GAT_OUT);
   G_2008GAT : Nor_gate port map( I1 => G_1908GAT_OUT, I2 => G_1955GAT_OUT, O 
                           => G_2008GAT_OUT);
   G_2007GAT : Nor_gate port map( I1 => G_1951GAT_OUT, I2 => G_1831GAT_OUT, O 
                           => G_2007GAT_OUT);
   G_2006GAT : Nor_gate port map( I1 => G_1905GAT_OUT, I2 => G_1951GAT_OUT, O 
                           => G_2006GAT_OUT);
   G_2005GAT : Nor_gate port map( I1 => G_1947GAT_OUT, I2 => G_1826GAT_OUT, O 
                           => G_2005GAT_OUT);
   G_2004GAT : Nor_gate port map( I1 => G_1902GAT_OUT, I2 => G_1947GAT_OUT, O 
                           => G_2004GAT_OUT);
   G_2001GAT : Nor_gate port map( I1 => G_1945GAT_OUT, I2 => G_1946GAT_OUT, O 
                           => G_2001GAT_OUT);
   G_2000GAT : Nor_gate port map( I1 => G_1941GAT_OUT, I2 => G_1891GAT_OUT, O 
                           => G_2000GAT_OUT);
   G_1999GAT : Nor_gate port map( I1 => G_1894GAT_OUT, I2 => G_1941GAT_OUT, O 
                           => G_1999GAT_OUT);
   G_1995GAT : Nor_gate port map( I1 => G_1938GAT_OUT, I2 => G_1886GAT_OUT, O 
                           => G_1995GAT_OUT);
   G_1991GAT : Nor_gate port map( I1 => G_1935GAT_OUT, I2 => G_1881GAT_OUT, O 
                           => G_1991GAT_OUT);
   G_1987GAT : Nor_gate port map( I1 => G_1932GAT_OUT, I2 => G_1876GAT_OUT, O 
                           => G_1987GAT_OUT);
   G_1983GAT : Nor_gate port map( I1 => G_1929GAT_OUT, I2 => G_1871GAT_OUT, O 
                           => G_1983GAT_OUT);
   G_1979GAT : Nor_gate port map( I1 => G_1926GAT_OUT, I2 => G_1866GAT_OUT, O 
                           => G_1979GAT_OUT);
   G_1975GAT : Nor_gate port map( I1 => G_1923GAT_OUT, I2 => G_1861GAT_OUT, O 
                           => G_1975GAT_OUT);
   G_1971GAT : Nor_gate port map( I1 => G_1920GAT_OUT, I2 => G_1856GAT_OUT, O 
                           => G_1971GAT_OUT);
   G_1967GAT : Nor_gate port map( I1 => G_1917GAT_OUT, I2 => G_1851GAT_OUT, O 
                           => G_1967GAT_OUT);
   G_1963GAT : Nor_gate port map( I1 => G_1914GAT_OUT, I2 => G_1846GAT_OUT, O 
                           => G_1963GAT_OUT);
   G_1959GAT : Nor_gate port map( I1 => G_1911GAT_OUT, I2 => G_1841GAT_OUT, O 
                           => G_1959GAT_OUT);
   G_1955GAT : Nor_gate port map( I1 => G_1908GAT_OUT, I2 => G_1836GAT_OUT, O 
                           => G_1955GAT_OUT);
   G_1951GAT : Nor_gate port map( I1 => G_1905GAT_OUT, I2 => G_1831GAT_OUT, O 
                           => G_1951GAT_OUT);
   G_1947GAT : Nor_gate port map( I1 => G_1902GAT_OUT, I2 => G_1826GAT_OUT, O 
                           => G_1947GAT_OUT);
   G_1946GAT : Nor_gate port map( I1 => G_1897GAT_OUT, I2 => G_1821GAT_OUT, O 
                           => G_1946GAT_OUT);
   G_1945GAT : Nor_gate port map( I1 => G_1269GAT_OUT, I2 => G_1897GAT_OUT, O 
                           => G_1945GAT_OUT);
   G_1941GAT : Nor_gate port map( I1 => G_1894GAT_OUT, I2 => G_1891GAT_OUT, O 
                           => G_1941GAT_OUT);
   G_1938GAT : Nor_gate port map( I1 => G_1889GAT_OUT, I2 => G_1890GAT_OUT, O 
                           => G_1938GAT_OUT);
   G_1935GAT : Nor_gate port map( I1 => G_1884GAT_OUT, I2 => G_1885GAT_OUT, O 
                           => G_1935GAT_OUT);
   G_1932GAT : Nor_gate port map( I1 => G_1879GAT_OUT, I2 => G_1880GAT_OUT, O 
                           => G_1932GAT_OUT);
   G_1929GAT : Nor_gate port map( I1 => G_1874GAT_OUT, I2 => G_1875GAT_OUT, O 
                           => G_1929GAT_OUT);
   G_1926GAT : Nor_gate port map( I1 => G_1869GAT_OUT, I2 => G_1870GAT_OUT, O 
                           => G_1926GAT_OUT);
   G_1923GAT : Nor_gate port map( I1 => G_1864GAT_OUT, I2 => G_1865GAT_OUT, O 
                           => G_1923GAT_OUT);
   G_1920GAT : Nor_gate port map( I1 => G_1859GAT_OUT, I2 => G_1860GAT_OUT, O 
                           => G_1920GAT_OUT);
   G_1917GAT : Nor_gate port map( I1 => G_1854GAT_OUT, I2 => G_1855GAT_OUT, O 
                           => G_1917GAT_OUT);
   G_1914GAT : Nor_gate port map( I1 => G_1849GAT_OUT, I2 => G_1850GAT_OUT, O 
                           => G_1914GAT_OUT);
   G_1911GAT : Nor_gate port map( I1 => G_1844GAT_OUT, I2 => G_1845GAT_OUT, O 
                           => G_1911GAT_OUT);
   G_1908GAT : Nor_gate port map( I1 => G_1839GAT_OUT, I2 => G_1840GAT_OUT, O 
                           => G_1908GAT_OUT);
   G_1905GAT : Nor_gate port map( I1 => G_1834GAT_OUT, I2 => G_1835GAT_OUT, O 
                           => G_1905GAT_OUT);
   G_1902GAT : Nor_gate port map( I1 => G_1829GAT_OUT, I2 => G_1830GAT_OUT, O 
                           => G_1902GAT_OUT);
   G_1897GAT : Nor_gate port map( I1 => G_1269GAT_OUT, I2 => G_1821GAT_OUT, O 
                           => G_1897GAT_OUT);
   G_1894GAT : Nor_gate port map( I1 => G_1819GAT_OUT, I2 => G_1820GAT_OUT, O 
                           => G_1894GAT_OUT);
   G_1891GAT : Nor_gate port map( I1 => G_1680GAT_OUT, I2 => G_1815GAT_OUT, O 
                           => G_1891GAT_OUT);
   G_1890GAT : Nor_gate port map( I1 => G_1815GAT_OUT, I2 => G_1173GAT_OUT, O 
                           => G_1890GAT_OUT);
   G_1889GAT : Nor_gate port map( I1 => G_1756GAT_OUT, I2 => G_1815GAT_OUT, O 
                           => G_1889GAT_OUT);
   G_1886GAT : Nor_gate port map( I1 => G_1676GAT_OUT, I2 => G_1811GAT_OUT, O 
                           => G_1886GAT_OUT);
   G_1885GAT : Nor_gate port map( I1 => G_1811GAT_OUT, I2 => G_1125GAT_OUT, O 
                           => G_1885GAT_OUT);
   G_1884GAT : Nor_gate port map( I1 => G_1753GAT_OUT, I2 => G_1811GAT_OUT, O 
                           => G_1884GAT_OUT);
   G_1881GAT : Nor_gate port map( I1 => G_1672GAT_OUT, I2 => G_1807GAT_OUT, O 
                           => G_1881GAT_OUT);
   G_1880GAT : Nor_gate port map( I1 => G_1807GAT_OUT, I2 => G_1077GAT_OUT, O 
                           => G_1880GAT_OUT);
   G_1879GAT : Nor_gate port map( I1 => G_1750GAT_OUT, I2 => G_1807GAT_OUT, O 
                           => G_1879GAT_OUT);
   G_1876GAT : Nor_gate port map( I1 => G_1668GAT_OUT, I2 => G_1803GAT_OUT, O 
                           => G_1876GAT_OUT);
   G_1875GAT : Nor_gate port map( I1 => G_1803GAT_OUT, I2 => G_1029GAT_OUT, O 
                           => G_1875GAT_OUT);
   G_1874GAT : Nor_gate port map( I1 => G_1747GAT_OUT, I2 => G_1803GAT_OUT, O 
                           => G_1874GAT_OUT);
   G_1871GAT : Nor_gate port map( I1 => G_1664GAT_OUT, I2 => G_1799GAT_OUT, O 
                           => G_1871GAT_OUT);
   G_1870GAT : Nor_gate port map( I1 => G_1799GAT_OUT, I2 => G_981GAT_OUT, O =>
                           G_1870GAT_OUT);
   G_1869GAT : Nor_gate port map( I1 => G_1744GAT_OUT, I2 => G_1799GAT_OUT, O 
                           => G_1869GAT_OUT);
   G_1866GAT : Nor_gate port map( I1 => G_1660GAT_OUT, I2 => G_1795GAT_OUT, O 
                           => G_1866GAT_OUT);
   G_1865GAT : Nor_gate port map( I1 => G_1795GAT_OUT, I2 => G_933GAT_OUT, O =>
                           G_1865GAT_OUT);
   G_1864GAT : Nor_gate port map( I1 => G_1741GAT_OUT, I2 => G_1795GAT_OUT, O 
                           => G_1864GAT_OUT);
   G_1861GAT : Nor_gate port map( I1 => G_1656GAT_OUT, I2 => G_1791GAT_OUT, O 
                           => G_1861GAT_OUT);
   G_1860GAT : Nor_gate port map( I1 => G_1791GAT_OUT, I2 => G_885GAT_OUT, O =>
                           G_1860GAT_OUT);
   G_1859GAT : Nor_gate port map( I1 => G_1738GAT_OUT, I2 => G_1791GAT_OUT, O 
                           => G_1859GAT_OUT);
   G_1856GAT : Nor_gate port map( I1 => G_1652GAT_OUT, I2 => G_1787GAT_OUT, O 
                           => G_1856GAT_OUT);
   G_1855GAT : Nor_gate port map( I1 => G_1787GAT_OUT, I2 => G_837GAT_OUT, O =>
                           G_1855GAT_OUT);
   G_1854GAT : Nor_gate port map( I1 => G_1735GAT_OUT, I2 => G_1787GAT_OUT, O 
                           => G_1854GAT_OUT);
   G_1851GAT : Nor_gate port map( I1 => G_1648GAT_OUT, I2 => G_1783GAT_OUT, O 
                           => G_1851GAT_OUT);
   G_1850GAT : Nor_gate port map( I1 => G_1783GAT_OUT, I2 => G_789GAT_OUT, O =>
                           G_1850GAT_OUT);
   G_1849GAT : Nor_gate port map( I1 => G_1732GAT_OUT, I2 => G_1783GAT_OUT, O 
                           => G_1849GAT_OUT);
   G_1846GAT : Nor_gate port map( I1 => G_1644GAT_OUT, I2 => G_1779GAT_OUT, O 
                           => G_1846GAT_OUT);
   G_1845GAT : Nor_gate port map( I1 => G_1779GAT_OUT, I2 => G_741GAT_OUT, O =>
                           G_1845GAT_OUT);
   G_1844GAT : Nor_gate port map( I1 => G_1729GAT_OUT, I2 => G_1779GAT_OUT, O 
                           => G_1844GAT_OUT);
   G_1841GAT : Nor_gate port map( I1 => G_1640GAT_OUT, I2 => G_1775GAT_OUT, O 
                           => G_1841GAT_OUT);
   G_1840GAT : Nor_gate port map( I1 => G_1775GAT_OUT, I2 => G_693GAT_OUT, O =>
                           G_1840GAT_OUT);
   G_1839GAT : Nor_gate port map( I1 => G_1726GAT_OUT, I2 => G_1775GAT_OUT, O 
                           => G_1839GAT_OUT);
   G_1836GAT : Nor_gate port map( I1 => G_1636GAT_OUT, I2 => G_1771GAT_OUT, O 
                           => G_1836GAT_OUT);
   G_1835GAT : Nor_gate port map( I1 => G_1771GAT_OUT, I2 => G_645GAT_OUT, O =>
                           G_1835GAT_OUT);
   G_1834GAT : Nor_gate port map( I1 => G_1723GAT_OUT, I2 => G_1771GAT_OUT, O 
                           => G_1834GAT_OUT);
   G_1831GAT : Nor_gate port map( I1 => G_1632GAT_OUT, I2 => G_1767GAT_OUT, O 
                           => G_1831GAT_OUT);
   G_1830GAT : Nor_gate port map( I1 => G_1767GAT_OUT, I2 => G_597GAT_OUT, O =>
                           G_1830GAT_OUT);
   G_1829GAT : Nor_gate port map( I1 => G_1720GAT_OUT, I2 => G_1767GAT_OUT, O 
                           => G_1829GAT_OUT);
   G_1826GAT : Nor_gate port map( I1 => G_1628GAT_OUT, I2 => G_1763GAT_OUT, O 
                           => G_1826GAT_OUT);
   G_1825GAT : Nor_gate port map( I1 => G_1763GAT_OUT, I2 => G_549GAT_OUT, O =>
                           G_1825GAT_OUT);
   G_1824GAT : Nor_gate port map( I1 => G_1717GAT_OUT, I2 => G_1763GAT_OUT, O 
                           => G_1824GAT_OUT);
   G_1821GAT : Nor_gate port map( I1 => G_1624GAT_OUT, I2 => G_1759GAT_OUT, O 
                           => G_1821GAT_OUT);
   G_1820GAT : Nor_gate port map( I1 => G_1759GAT_OUT, I2 => G_1221GAT_OUT, O 
                           => G_1820GAT_OUT);
   G_1819GAT : Nor_gate port map( I1 => G_1714GAT_OUT, I2 => G_1759GAT_OUT, O 
                           => G_1819GAT_OUT);
   G_1815GAT : Nor_gate port map( I1 => G_1756GAT_OUT, I2 => G_1173GAT_OUT, O 
                           => G_1815GAT_OUT);
   G_1811GAT : Nor_gate port map( I1 => G_1753GAT_OUT, I2 => G_1125GAT_OUT, O 
                           => G_1811GAT_OUT);
   G_1807GAT : Nor_gate port map( I1 => G_1750GAT_OUT, I2 => G_1077GAT_OUT, O 
                           => G_1807GAT_OUT);
   G_1803GAT : Nor_gate port map( I1 => G_1747GAT_OUT, I2 => G_1029GAT_OUT, O 
                           => G_1803GAT_OUT);
   G_1799GAT : Nor_gate port map( I1 => G_1744GAT_OUT, I2 => G_981GAT_OUT, O =>
                           G_1799GAT_OUT);
   G_1795GAT : Nor_gate port map( I1 => G_1741GAT_OUT, I2 => G_933GAT_OUT, O =>
                           G_1795GAT_OUT);
   G_1791GAT : Nor_gate port map( I1 => G_1738GAT_OUT, I2 => G_885GAT_OUT, O =>
                           G_1791GAT_OUT);
   G_1787GAT : Nor_gate port map( I1 => G_1735GAT_OUT, I2 => G_837GAT_OUT, O =>
                           G_1787GAT_OUT);
   G_1783GAT : Nor_gate port map( I1 => G_1732GAT_OUT, I2 => G_789GAT_OUT, O =>
                           G_1783GAT_OUT);
   G_1779GAT : Nor_gate port map( I1 => G_1729GAT_OUT, I2 => G_741GAT_OUT, O =>
                           G_1779GAT_OUT);
   G_1775GAT : Nor_gate port map( I1 => G_1726GAT_OUT, I2 => G_693GAT_OUT, O =>
                           G_1775GAT_OUT);
   G_1771GAT : Nor_gate port map( I1 => G_1723GAT_OUT, I2 => G_645GAT_OUT, O =>
                           G_1771GAT_OUT);
   G_1767GAT : Nor_gate port map( I1 => G_1720GAT_OUT, I2 => G_597GAT_OUT, O =>
                           G_1767GAT_OUT);
   G_1763GAT : Nor_gate port map( I1 => G_1717GAT_OUT, I2 => G_549GAT_OUT, O =>
                           G_1763GAT_OUT);
   G_1759GAT : Nor_gate port map( I1 => G_1714GAT_OUT, I2 => G_1221GAT_OUT, O 
                           => G_1759GAT_OUT);
   G_1756GAT : Nor_gate port map( I1 => G_1712GAT_OUT, I2 => G_1713GAT_OUT, O 
                           => G_1756GAT_OUT);
   G_1753GAT : Nor_gate port map( I1 => G_1710GAT_OUT, I2 => G_1711GAT_OUT, O 
                           => G_1753GAT_OUT);
   G_1750GAT : Nor_gate port map( I1 => G_1708GAT_OUT, I2 => G_1709GAT_OUT, O 
                           => G_1750GAT_OUT);
   G_1747GAT : Nor_gate port map( I1 => G_1706GAT_OUT, I2 => G_1707GAT_OUT, O 
                           => G_1747GAT_OUT);
   G_1744GAT : Nor_gate port map( I1 => G_1704GAT_OUT, I2 => G_1705GAT_OUT, O 
                           => G_1744GAT_OUT);
   G_1741GAT : Nor_gate port map( I1 => G_1702GAT_OUT, I2 => G_1703GAT_OUT, O 
                           => G_1741GAT_OUT);
   G_1738GAT : Nor_gate port map( I1 => G_1700GAT_OUT, I2 => G_1701GAT_OUT, O 
                           => G_1738GAT_OUT);
   G_1735GAT : Nor_gate port map( I1 => G_1698GAT_OUT, I2 => G_1699GAT_OUT, O 
                           => G_1735GAT_OUT);
   G_1732GAT : Nor_gate port map( I1 => G_1696GAT_OUT, I2 => G_1697GAT_OUT, O 
                           => G_1732GAT_OUT);
   G_1729GAT : Nor_gate port map( I1 => G_1694GAT_OUT, I2 => G_1695GAT_OUT, O 
                           => G_1729GAT_OUT);
   G_1726GAT : Nor_gate port map( I1 => G_1692GAT_OUT, I2 => G_1693GAT_OUT, O 
                           => G_1726GAT_OUT);
   G_1723GAT : Nor_gate port map( I1 => G_1690GAT_OUT, I2 => G_1691GAT_OUT, O 
                           => G_1723GAT_OUT);
   G_1720GAT : Nor_gate port map( I1 => G_1688GAT_OUT, I2 => G_1689GAT_OUT, O 
                           => G_1720GAT_OUT);
   G_1717GAT : Nor_gate port map( I1 => G_1686GAT_OUT, I2 => G_1687GAT_OUT, O 
                           => G_1717GAT_OUT);
   G_1714GAT : Nor_gate port map( I1 => G_1684GAT_OUT, I2 => G_1685GAT_OUT, O 
                           => G_1714GAT_OUT);
   G_1713GAT : Nor_gate port map( I1 => G_1680GAT_OUT, I2 => G_1573GAT_OUT, O 
                           => G_1713GAT_OUT);
   G_1712GAT : Nor_gate port map( I1 => G_1621GAT_OUT, I2 => G_1680GAT_OUT, O 
                           => G_1712GAT_OUT);
   G_1711GAT : Nor_gate port map( I1 => G_1676GAT_OUT, I2 => G_1568GAT_OUT, O 
                           => G_1711GAT_OUT);
   G_1710GAT : Nor_gate port map( I1 => G_1618GAT_OUT, I2 => G_1676GAT_OUT, O 
                           => G_1710GAT_OUT);
   G_1709GAT : Nor_gate port map( I1 => G_1672GAT_OUT, I2 => G_1563GAT_OUT, O 
                           => G_1709GAT_OUT);
   G_1708GAT : Nor_gate port map( I1 => G_1615GAT_OUT, I2 => G_1672GAT_OUT, O 
                           => G_1708GAT_OUT);
   G_1707GAT : Nor_gate port map( I1 => G_1668GAT_OUT, I2 => G_1558GAT_OUT, O 
                           => G_1707GAT_OUT);
   G_1706GAT : Nor_gate port map( I1 => G_1612GAT_OUT, I2 => G_1668GAT_OUT, O 
                           => G_1706GAT_OUT);
   G_1705GAT : Nor_gate port map( I1 => G_1664GAT_OUT, I2 => G_1553GAT_OUT, O 
                           => G_1705GAT_OUT);
   G_1704GAT : Nor_gate port map( I1 => G_1609GAT_OUT, I2 => G_1664GAT_OUT, O 
                           => G_1704GAT_OUT);
   G_1703GAT : Nor_gate port map( I1 => G_1660GAT_OUT, I2 => G_1548GAT_OUT, O 
                           => G_1703GAT_OUT);
   G_1702GAT : Nor_gate port map( I1 => G_1606GAT_OUT, I2 => G_1660GAT_OUT, O 
                           => G_1702GAT_OUT);
   G_1701GAT : Nor_gate port map( I1 => G_1656GAT_OUT, I2 => G_1543GAT_OUT, O 
                           => G_1701GAT_OUT);
   G_1700GAT : Nor_gate port map( I1 => G_1603GAT_OUT, I2 => G_1656GAT_OUT, O 
                           => G_1700GAT_OUT);
   G_1699GAT : Nor_gate port map( I1 => G_1652GAT_OUT, I2 => G_1538GAT_OUT, O 
                           => G_1699GAT_OUT);
   G_1698GAT : Nor_gate port map( I1 => G_1600GAT_OUT, I2 => G_1652GAT_OUT, O 
                           => G_1698GAT_OUT);
   G_1697GAT : Nor_gate port map( I1 => G_1648GAT_OUT, I2 => G_1533GAT_OUT, O 
                           => G_1697GAT_OUT);
   G_1696GAT : Nor_gate port map( I1 => G_1597GAT_OUT, I2 => G_1648GAT_OUT, O 
                           => G_1696GAT_OUT);
   G_1695GAT : Nor_gate port map( I1 => G_1644GAT_OUT, I2 => G_1528GAT_OUT, O 
                           => G_1695GAT_OUT);
   G_1694GAT : Nor_gate port map( I1 => G_1594GAT_OUT, I2 => G_1644GAT_OUT, O 
                           => G_1694GAT_OUT);
   G_1693GAT : Nor_gate port map( I1 => G_1640GAT_OUT, I2 => G_1523GAT_OUT, O 
                           => G_1693GAT_OUT);
   G_1692GAT : Nor_gate port map( I1 => G_1591GAT_OUT, I2 => G_1640GAT_OUT, O 
                           => G_1692GAT_OUT);
   G_1691GAT : Nor_gate port map( I1 => G_1636GAT_OUT, I2 => G_1518GAT_OUT, O 
                           => G_1691GAT_OUT);
   G_1690GAT : Nor_gate port map( I1 => G_1588GAT_OUT, I2 => G_1636GAT_OUT, O 
                           => G_1690GAT_OUT);
   G_1689GAT : Nor_gate port map( I1 => G_1632GAT_OUT, I2 => G_1513GAT_OUT, O 
                           => G_1689GAT_OUT);
   G_1688GAT : Nor_gate port map( I1 => G_1585GAT_OUT, I2 => G_1632GAT_OUT, O 
                           => G_1688GAT_OUT);
   G_1687GAT : Nor_gate port map( I1 => G_1628GAT_OUT, I2 => G_1508GAT_OUT, O 
                           => G_1687GAT_OUT);
   G_1686GAT : Nor_gate port map( I1 => G_1582GAT_OUT, I2 => G_1628GAT_OUT, O 
                           => G_1686GAT_OUT);
   G_1685GAT : Nor_gate port map( I1 => G_1624GAT_OUT, I2 => G_1578GAT_OUT, O 
                           => G_1685GAT_OUT);
   G_1684GAT : Nor_gate port map( I1 => G_1266GAT_OUT, I2 => G_1624GAT_OUT, O 
                           => G_1684GAT_OUT);
   G_1680GAT : Nor_gate port map( I1 => G_1621GAT_OUT, I2 => G_1573GAT_OUT, O 
                           => G_1680GAT_OUT);
   G_1676GAT : Nor_gate port map( I1 => G_1618GAT_OUT, I2 => G_1568GAT_OUT, O 
                           => G_1676GAT_OUT);
   G_1672GAT : Nor_gate port map( I1 => G_1615GAT_OUT, I2 => G_1563GAT_OUT, O 
                           => G_1672GAT_OUT);
   G_1668GAT : Nor_gate port map( I1 => G_1612GAT_OUT, I2 => G_1558GAT_OUT, O 
                           => G_1668GAT_OUT);
   G_1664GAT : Nor_gate port map( I1 => G_1609GAT_OUT, I2 => G_1553GAT_OUT, O 
                           => G_1664GAT_OUT);
   G_1660GAT : Nor_gate port map( I1 => G_1606GAT_OUT, I2 => G_1548GAT_OUT, O 
                           => G_1660GAT_OUT);
   G_1656GAT : Nor_gate port map( I1 => G_1603GAT_OUT, I2 => G_1543GAT_OUT, O 
                           => G_1656GAT_OUT);
   G_1652GAT : Nor_gate port map( I1 => G_1600GAT_OUT, I2 => G_1538GAT_OUT, O 
                           => G_1652GAT_OUT);
   G_1648GAT : Nor_gate port map( I1 => G_1597GAT_OUT, I2 => G_1533GAT_OUT, O 
                           => G_1648GAT_OUT);
   G_1644GAT : Nor_gate port map( I1 => G_1594GAT_OUT, I2 => G_1528GAT_OUT, O 
                           => G_1644GAT_OUT);
   G_1640GAT : Nor_gate port map( I1 => G_1591GAT_OUT, I2 => G_1523GAT_OUT, O 
                           => G_1640GAT_OUT);
   G_1636GAT : Nor_gate port map( I1 => G_1588GAT_OUT, I2 => G_1518GAT_OUT, O 
                           => G_1636GAT_OUT);
   G_1632GAT : Nor_gate port map( I1 => G_1585GAT_OUT, I2 => G_1513GAT_OUT, O 
                           => G_1632GAT_OUT);
   G_1628GAT : Nor_gate port map( I1 => G_1582GAT_OUT, I2 => G_1508GAT_OUT, O 
                           => G_1628GAT_OUT);
   G_1624GAT : Nor_gate port map( I1 => G_1266GAT_OUT, I2 => G_1578GAT_OUT, O 
                           => G_1624GAT_OUT);
   G_1621GAT : Nor_gate port map( I1 => G_1576GAT_OUT, I2 => G_1577GAT_OUT, O 
                           => G_1621GAT_OUT);
   G_1618GAT : Nor_gate port map( I1 => G_1571GAT_OUT, I2 => G_1572GAT_OUT, O 
                           => G_1618GAT_OUT);
   G_1615GAT : Nor_gate port map( I1 => G_1566GAT_OUT, I2 => G_1567GAT_OUT, O 
                           => G_1615GAT_OUT);
   G_1612GAT : Nor_gate port map( I1 => G_1561GAT_OUT, I2 => G_1562GAT_OUT, O 
                           => G_1612GAT_OUT);
   G_1609GAT : Nor_gate port map( I1 => G_1556GAT_OUT, I2 => G_1557GAT_OUT, O 
                           => G_1609GAT_OUT);
   G_1606GAT : Nor_gate port map( I1 => G_1551GAT_OUT, I2 => G_1552GAT_OUT, O 
                           => G_1606GAT_OUT);
   G_1603GAT : Nor_gate port map( I1 => G_1546GAT_OUT, I2 => G_1547GAT_OUT, O 
                           => G_1603GAT_OUT);
   G_1600GAT : Nor_gate port map( I1 => G_1541GAT_OUT, I2 => G_1542GAT_OUT, O 
                           => G_1600GAT_OUT);
   G_1597GAT : Nor_gate port map( I1 => G_1536GAT_OUT, I2 => G_1537GAT_OUT, O 
                           => G_1597GAT_OUT);
   G_1594GAT : Nor_gate port map( I1 => G_1531GAT_OUT, I2 => G_1532GAT_OUT, O 
                           => G_1594GAT_OUT);
   G_1591GAT : Nor_gate port map( I1 => G_1526GAT_OUT, I2 => G_1527GAT_OUT, O 
                           => G_1591GAT_OUT);
   G_1588GAT : Nor_gate port map( I1 => G_1521GAT_OUT, I2 => G_1522GAT_OUT, O 
                           => G_1588GAT_OUT);
   G_1585GAT : Nor_gate port map( I1 => G_1516GAT_OUT, I2 => G_1517GAT_OUT, O 
                           => G_1585GAT_OUT);
   G_1582GAT : Nor_gate port map( I1 => G_1511GAT_OUT, I2 => G_1512GAT_OUT, O 
                           => G_1582GAT_OUT);
   G_1578GAT : Nor_gate port map( I1 => G_1367GAT_OUT, I2 => G_1502GAT_OUT, O 
                           => G_1578GAT_OUT);
   G_1577GAT : Nor_gate port map( I1 => G_1502GAT_OUT, I2 => G_1218GAT_OUT, O 
                           => G_1577GAT_OUT);
   G_1576GAT : Nor_gate port map( I1 => G_1443GAT_OUT, I2 => G_1502GAT_OUT, O 
                           => G_1576GAT_OUT);
   G_1573GAT : Nor_gate port map( I1 => G_1363GAT_OUT, I2 => G_1498GAT_OUT, O 
                           => G_1573GAT_OUT);
   G_1572GAT : Nor_gate port map( I1 => G_1498GAT_OUT, I2 => G_1170GAT_OUT, O 
                           => G_1572GAT_OUT);
   G_1571GAT : Nor_gate port map( I1 => G_1440GAT_OUT, I2 => G_1498GAT_OUT, O 
                           => G_1571GAT_OUT);
   G_1568GAT : Nor_gate port map( I1 => G_1359GAT_OUT, I2 => G_1494GAT_OUT, O 
                           => G_1568GAT_OUT);
   G_1567GAT : Nor_gate port map( I1 => G_1494GAT_OUT, I2 => G_1122GAT_OUT, O 
                           => G_1567GAT_OUT);
   G_1566GAT : Nor_gate port map( I1 => G_1437GAT_OUT, I2 => G_1494GAT_OUT, O 
                           => G_1566GAT_OUT);
   G_1563GAT : Nor_gate port map( I1 => G_1355GAT_OUT, I2 => G_1490GAT_OUT, O 
                           => G_1563GAT_OUT);
   G_1562GAT : Nor_gate port map( I1 => G_1490GAT_OUT, I2 => G_1074GAT_OUT, O 
                           => G_1562GAT_OUT);
   G_1561GAT : Nor_gate port map( I1 => G_1434GAT_OUT, I2 => G_1490GAT_OUT, O 
                           => G_1561GAT_OUT);
   G_1558GAT : Nor_gate port map( I1 => G_1351GAT_OUT, I2 => G_1486GAT_OUT, O 
                           => G_1558GAT_OUT);
   G_1557GAT : Nor_gate port map( I1 => G_1486GAT_OUT, I2 => G_1026GAT_OUT, O 
                           => G_1557GAT_OUT);
   G_1556GAT : Nor_gate port map( I1 => G_1431GAT_OUT, I2 => G_1486GAT_OUT, O 
                           => G_1556GAT_OUT);
   G_1553GAT : Nor_gate port map( I1 => G_1347GAT_OUT, I2 => G_1482GAT_OUT, O 
                           => G_1553GAT_OUT);
   G_1552GAT : Nor_gate port map( I1 => G_1482GAT_OUT, I2 => G_978GAT_OUT, O =>
                           G_1552GAT_OUT);
   G_1551GAT : Nor_gate port map( I1 => G_1428GAT_OUT, I2 => G_1482GAT_OUT, O 
                           => G_1551GAT_OUT);
   G_1548GAT : Nor_gate port map( I1 => G_1343GAT_OUT, I2 => G_1478GAT_OUT, O 
                           => G_1548GAT_OUT);
   G_1547GAT : Nor_gate port map( I1 => G_1478GAT_OUT, I2 => G_930GAT_OUT, O =>
                           G_1547GAT_OUT);
   G_1546GAT : Nor_gate port map( I1 => G_1425GAT_OUT, I2 => G_1478GAT_OUT, O 
                           => G_1546GAT_OUT);
   G_1543GAT : Nor_gate port map( I1 => G_1339GAT_OUT, I2 => G_1474GAT_OUT, O 
                           => G_1543GAT_OUT);
   G_1542GAT : Nor_gate port map( I1 => G_1474GAT_OUT, I2 => G_882GAT_OUT, O =>
                           G_1542GAT_OUT);
   G_1541GAT : Nor_gate port map( I1 => G_1422GAT_OUT, I2 => G_1474GAT_OUT, O 
                           => G_1541GAT_OUT);
   G_1538GAT : Nor_gate port map( I1 => G_1335GAT_OUT, I2 => G_1470GAT_OUT, O 
                           => G_1538GAT_OUT);
   G_1537GAT : Nor_gate port map( I1 => G_1470GAT_OUT, I2 => G_834GAT_OUT, O =>
                           G_1537GAT_OUT);
   G_1536GAT : Nor_gate port map( I1 => G_1419GAT_OUT, I2 => G_1470GAT_OUT, O 
                           => G_1536GAT_OUT);
   G_1533GAT : Nor_gate port map( I1 => G_1331GAT_OUT, I2 => G_1466GAT_OUT, O 
                           => G_1533GAT_OUT);
   G_1532GAT : Nor_gate port map( I1 => G_1466GAT_OUT, I2 => G_786GAT_OUT, O =>
                           G_1532GAT_OUT);
   G_1531GAT : Nor_gate port map( I1 => G_1416GAT_OUT, I2 => G_1466GAT_OUT, O 
                           => G_1531GAT_OUT);
   G_1528GAT : Nor_gate port map( I1 => G_1327GAT_OUT, I2 => G_1462GAT_OUT, O 
                           => G_1528GAT_OUT);
   G_1527GAT : Nor_gate port map( I1 => G_1462GAT_OUT, I2 => G_738GAT_OUT, O =>
                           G_1527GAT_OUT);
   G_1526GAT : Nor_gate port map( I1 => G_1413GAT_OUT, I2 => G_1462GAT_OUT, O 
                           => G_1526GAT_OUT);
   G_1523GAT : Nor_gate port map( I1 => G_1323GAT_OUT, I2 => G_1458GAT_OUT, O 
                           => G_1523GAT_OUT);
   G_1522GAT : Nor_gate port map( I1 => G_1458GAT_OUT, I2 => G_690GAT_OUT, O =>
                           G_1522GAT_OUT);
   G_1521GAT : Nor_gate port map( I1 => G_1410GAT_OUT, I2 => G_1458GAT_OUT, O 
                           => G_1521GAT_OUT);
   G_1518GAT : Nor_gate port map( I1 => G_1319GAT_OUT, I2 => G_1454GAT_OUT, O 
                           => G_1518GAT_OUT);
   G_1517GAT : Nor_gate port map( I1 => G_1454GAT_OUT, I2 => G_642GAT_OUT, O =>
                           G_1517GAT_OUT);
   G_1516GAT : Nor_gate port map( I1 => G_1407GAT_OUT, I2 => G_1454GAT_OUT, O 
                           => G_1516GAT_OUT);
   G_1513GAT : Nor_gate port map( I1 => G_1315GAT_OUT, I2 => G_1450GAT_OUT, O 
                           => G_1513GAT_OUT);
   G_1512GAT : Nor_gate port map( I1 => G_1450GAT_OUT, I2 => G_594GAT_OUT, O =>
                           G_1512GAT_OUT);
   G_1511GAT : Nor_gate port map( I1 => G_1404GAT_OUT, I2 => G_1450GAT_OUT, O 
                           => G_1511GAT_OUT);
   G_1508GAT : Nor_gate port map( I1 => G_1311GAT_OUT, I2 => G_1446GAT_OUT, O 
                           => G_1508GAT_OUT);
   G_1507GAT : Nor_gate port map( I1 => G_1446GAT_OUT, I2 => G_546GAT_OUT, O =>
                           G_1507GAT_OUT);
   G_1506GAT : Nor_gate port map( I1 => G_1401GAT_OUT, I2 => G_1446GAT_OUT, O 
                           => G_1506GAT_OUT);
   G_1502GAT : Nor_gate port map( I1 => G_1443GAT_OUT, I2 => G_1218GAT_OUT, O 
                           => G_1502GAT_OUT);
   G_1498GAT : Nor_gate port map( I1 => G_1440GAT_OUT, I2 => G_1170GAT_OUT, O 
                           => G_1498GAT_OUT);
   G_1494GAT : Nor_gate port map( I1 => G_1437GAT_OUT, I2 => G_1122GAT_OUT, O 
                           => G_1494GAT_OUT);
   G_1490GAT : Nor_gate port map( I1 => G_1434GAT_OUT, I2 => G_1074GAT_OUT, O 
                           => G_1490GAT_OUT);
   G_1486GAT : Nor_gate port map( I1 => G_1431GAT_OUT, I2 => G_1026GAT_OUT, O 
                           => G_1486GAT_OUT);
   G_1482GAT : Nor_gate port map( I1 => G_1428GAT_OUT, I2 => G_978GAT_OUT, O =>
                           G_1482GAT_OUT);
   G_1478GAT : Nor_gate port map( I1 => G_1425GAT_OUT, I2 => G_930GAT_OUT, O =>
                           G_1478GAT_OUT);
   G_1474GAT : Nor_gate port map( I1 => G_1422GAT_OUT, I2 => G_882GAT_OUT, O =>
                           G_1474GAT_OUT);
   G_1470GAT : Nor_gate port map( I1 => G_1419GAT_OUT, I2 => G_834GAT_OUT, O =>
                           G_1470GAT_OUT);
   G_1466GAT : Nor_gate port map( I1 => G_1416GAT_OUT, I2 => G_786GAT_OUT, O =>
                           G_1466GAT_OUT);
   G_1462GAT : Nor_gate port map( I1 => G_1413GAT_OUT, I2 => G_738GAT_OUT, O =>
                           G_1462GAT_OUT);
   G_1458GAT : Nor_gate port map( I1 => G_1410GAT_OUT, I2 => G_690GAT_OUT, O =>
                           G_1458GAT_OUT);
   G_1454GAT : Nor_gate port map( I1 => G_1407GAT_OUT, I2 => G_642GAT_OUT, O =>
                           G_1454GAT_OUT);
   G_1450GAT : Nor_gate port map( I1 => G_1404GAT_OUT, I2 => G_594GAT_OUT, O =>
                           G_1450GAT_OUT);
   G_1446GAT : Nor_gate port map( I1 => G_1401GAT_OUT, I2 => G_546GAT_OUT, O =>
                           G_1446GAT_OUT);
   G_1443GAT : Nor_gate port map( I1 => G_1399GAT_OUT, I2 => G_1400GAT_OUT, O 
                           => G_1443GAT_OUT);
   G_1440GAT : Nor_gate port map( I1 => G_1397GAT_OUT, I2 => G_1398GAT_OUT, O 
                           => G_1440GAT_OUT);
   G_1437GAT : Nor_gate port map( I1 => G_1395GAT_OUT, I2 => G_1396GAT_OUT, O 
                           => G_1437GAT_OUT);
   G_1434GAT : Nor_gate port map( I1 => G_1393GAT_OUT, I2 => G_1394GAT_OUT, O 
                           => G_1434GAT_OUT);
   G_1431GAT : Nor_gate port map( I1 => G_1391GAT_OUT, I2 => G_1392GAT_OUT, O 
                           => G_1431GAT_OUT);
   G_1428GAT : Nor_gate port map( I1 => G_1389GAT_OUT, I2 => G_1390GAT_OUT, O 
                           => G_1428GAT_OUT);
   G_1425GAT : Nor_gate port map( I1 => G_1387GAT_OUT, I2 => G_1388GAT_OUT, O 
                           => G_1425GAT_OUT);
   G_1422GAT : Nor_gate port map( I1 => G_1385GAT_OUT, I2 => G_1386GAT_OUT, O 
                           => G_1422GAT_OUT);
   G_1419GAT : Nor_gate port map( I1 => G_1383GAT_OUT, I2 => G_1384GAT_OUT, O 
                           => G_1419GAT_OUT);
   G_1416GAT : Nor_gate port map( I1 => G_1381GAT_OUT, I2 => G_1382GAT_OUT, O 
                           => G_1416GAT_OUT);
   G_1413GAT : Nor_gate port map( I1 => G_1379GAT_OUT, I2 => G_1380GAT_OUT, O 
                           => G_1413GAT_OUT);
   G_1410GAT : Nor_gate port map( I1 => G_1377GAT_OUT, I2 => G_1378GAT_OUT, O 
                           => G_1410GAT_OUT);
   G_1407GAT : Nor_gate port map( I1 => G_1375GAT_OUT, I2 => G_1376GAT_OUT, O 
                           => G_1407GAT_OUT);
   G_1404GAT : Nor_gate port map( I1 => G_1373GAT_OUT, I2 => G_1374GAT_OUT, O 
                           => G_1404GAT_OUT);
   G_1401GAT : Nor_gate port map( I1 => G_1371GAT_OUT, I2 => G_1372GAT_OUT, O 
                           => G_1401GAT_OUT);
   G_1400GAT : Inv_gate port map( I1 => G_1367GAT_OUT, O => G_1400GAT_OUT);
   G_1399GAT : Nor_gate port map( I1 => G_1263GAT_OUT, I2 => G_1367GAT_OUT, O 
                           => G_1399GAT_OUT);
   G_1398GAT : Inv_gate port map( I1 => G_1363GAT_OUT, O => G_1398GAT_OUT);
   G_1397GAT : Nor_gate port map( I1 => G_1215GAT_OUT, I2 => G_1363GAT_OUT, O 
                           => G_1397GAT_OUT);
   G_1396GAT : Inv_gate port map( I1 => G_1359GAT_OUT, O => G_1396GAT_OUT);
   G_1395GAT : Nor_gate port map( I1 => G_1167GAT_OUT, I2 => G_1359GAT_OUT, O 
                           => G_1395GAT_OUT);
   G_1394GAT : Inv_gate port map( I1 => G_1355GAT_OUT, O => G_1394GAT_OUT);
   G_1393GAT : Nor_gate port map( I1 => G_1119GAT_OUT, I2 => G_1355GAT_OUT, O 
                           => G_1393GAT_OUT);
   G_1392GAT : Inv_gate port map( I1 => G_1351GAT_OUT, O => G_1392GAT_OUT);
   G_1391GAT : Nor_gate port map( I1 => G_1071GAT_OUT, I2 => G_1351GAT_OUT, O 
                           => G_1391GAT_OUT);
   G_1390GAT : Inv_gate port map( I1 => G_1347GAT_OUT, O => G_1390GAT_OUT);
   G_1389GAT : Nor_gate port map( I1 => G_1023GAT_OUT, I2 => G_1347GAT_OUT, O 
                           => G_1389GAT_OUT);
   G_1388GAT : Inv_gate port map( I1 => G_1343GAT_OUT, O => G_1388GAT_OUT);
   G_1387GAT : Nor_gate port map( I1 => G_975GAT_OUT, I2 => G_1343GAT_OUT, O =>
                           G_1387GAT_OUT);
   G_1386GAT : Inv_gate port map( I1 => G_1339GAT_OUT, O => G_1386GAT_OUT);
   G_1385GAT : Nor_gate port map( I1 => G_927GAT_OUT, I2 => G_1339GAT_OUT, O =>
                           G_1385GAT_OUT);
   G_1384GAT : Inv_gate port map( I1 => G_1335GAT_OUT, O => G_1384GAT_OUT);
   G_1383GAT : Nor_gate port map( I1 => G_879GAT_OUT, I2 => G_1335GAT_OUT, O =>
                           G_1383GAT_OUT);
   G_1382GAT : Inv_gate port map( I1 => G_1331GAT_OUT, O => G_1382GAT_OUT);
   G_1381GAT : Nor_gate port map( I1 => G_831GAT_OUT, I2 => G_1331GAT_OUT, O =>
                           G_1381GAT_OUT);
   G_1380GAT : Inv_gate port map( I1 => G_1327GAT_OUT, O => G_1380GAT_OUT);
   G_1379GAT : Nor_gate port map( I1 => G_783GAT_OUT, I2 => G_1327GAT_OUT, O =>
                           G_1379GAT_OUT);
   G_1378GAT : Inv_gate port map( I1 => G_1323GAT_OUT, O => G_1378GAT_OUT);
   G_1377GAT : Nor_gate port map( I1 => G_735GAT_OUT, I2 => G_1323GAT_OUT, O =>
                           G_1377GAT_OUT);
   G_1376GAT : Inv_gate port map( I1 => G_1319GAT_OUT, O => G_1376GAT_OUT);
   G_1375GAT : Nor_gate port map( I1 => G_687GAT_OUT, I2 => G_1319GAT_OUT, O =>
                           G_1375GAT_OUT);
   G_1374GAT : Inv_gate port map( I1 => G_1315GAT_OUT, O => G_1374GAT_OUT);
   G_1373GAT : Nor_gate port map( I1 => G_639GAT_OUT, I2 => G_1315GAT_OUT, O =>
                           G_1373GAT_OUT);
   G_1372GAT : Inv_gate port map( I1 => G_1311GAT_OUT, O => G_1372GAT_OUT);
   G_1371GAT : Nor_gate port map( I1 => G_591GAT_OUT, I2 => G_1311GAT_OUT, O =>
                           G_1371GAT_OUT);
   G_1367GAT : Inv_gate port map( I1 => G_1263GAT_OUT, O => G_1367GAT_OUT);
   G_1363GAT : Inv_gate port map( I1 => G_1215GAT_OUT, O => G_1363GAT_OUT);
   G_1359GAT : Inv_gate port map( I1 => G_1167GAT_OUT, O => G_1359GAT_OUT);
   G_1355GAT : Inv_gate port map( I1 => G_1119GAT_OUT, O => G_1355GAT_OUT);
   G_1351GAT : Inv_gate port map( I1 => G_1071GAT_OUT, O => G_1351GAT_OUT);
   G_1347GAT : Inv_gate port map( I1 => G_1023GAT_OUT, O => G_1347GAT_OUT);
   G_1343GAT : Inv_gate port map( I1 => G_975GAT_OUT, O => G_1343GAT_OUT);
   G_1339GAT : Inv_gate port map( I1 => G_927GAT_OUT, O => G_1339GAT_OUT);
   G_1335GAT : Inv_gate port map( I1 => G_879GAT_OUT, O => G_1335GAT_OUT);
   G_1331GAT : Inv_gate port map( I1 => G_831GAT_OUT, O => G_1331GAT_OUT);
   G_1327GAT : Inv_gate port map( I1 => G_783GAT_OUT, O => G_1327GAT_OUT);
   G_1323GAT : Inv_gate port map( I1 => G_735GAT_OUT, O => G_1323GAT_OUT);
   G_1319GAT : Inv_gate port map( I1 => G_687GAT_OUT, O => G_1319GAT_OUT);
   G_1315GAT : Inv_gate port map( I1 => G_639GAT_OUT, O => G_1315GAT_OUT);
   G_1311GAT : Inv_gate port map( I1 => G_591GAT_OUT, O => G_1311GAT_OUT);
   G_1308GAT : And_gate port map( I1 => G_256GAT, I2 => G_528GAT, O => 
                           G_1308GAT_OUT);
   G_1305GAT : And_gate port map( I1 => G_256GAT, I2 => G_511GAT, O => 
                           G_1305GAT_OUT);
   G_1302GAT : And_gate port map( I1 => G_256GAT, I2 => G_494GAT, O => 
                           G_1302GAT_OUT);
   G_1299GAT : And_gate port map( I1 => G_256GAT, I2 => G_477GAT, O => 
                           G_1299GAT_OUT);
   G_1296GAT : And_gate port map( I1 => G_256GAT, I2 => G_460GAT, O => 
                           G_1296GAT_OUT);
   G_1293GAT : And_gate port map( I1 => G_256GAT, I2 => G_443GAT, O => 
                           G_1293GAT_OUT);
   G_1290GAT : And_gate port map( I1 => G_256GAT, I2 => G_426GAT, O => 
                           G_1290GAT_OUT);
   G_1287GAT : And_gate port map( I1 => G_256GAT, I2 => G_409GAT, O => 
                           G_1287GAT_OUT);
   G_1284GAT : And_gate port map( I1 => G_256GAT, I2 => G_392GAT, O => 
                           G_1284GAT_OUT);
   G_1281GAT : And_gate port map( I1 => G_256GAT, I2 => G_375GAT, O => 
                           G_1281GAT_OUT);
   G_1278GAT : And_gate port map( I1 => G_256GAT, I2 => G_358GAT, O => 
                           G_1278GAT_OUT);
   G_1275GAT : And_gate port map( I1 => G_256GAT, I2 => G_341GAT, O => 
                           G_1275GAT_OUT);
   G_1272GAT : And_gate port map( I1 => G_256GAT, I2 => G_324GAT, O => 
                           G_1272GAT_OUT);
   G_1269GAT : And_gate port map( I1 => G_256GAT, I2 => G_307GAT, O => 
                           G_1269GAT_OUT);
   G_1266GAT : And_gate port map( I1 => G_256GAT, I2 => G_290GAT, O => 
                           G_1266GAT_OUT);
   G_1263GAT : And_gate port map( I1 => G_256GAT, I2 => G_273GAT, O => 
                           G_1263GAT_OUT);
   G_1260GAT : And_gate port map( I1 => G_239GAT, I2 => G_528GAT, O => 
                           G_1260GAT_OUT);
   G_1257GAT : And_gate port map( I1 => G_239GAT, I2 => G_511GAT, O => 
                           G_1257GAT_OUT);
   G_1254GAT : And_gate port map( I1 => G_239GAT, I2 => G_494GAT, O => 
                           G_1254GAT_OUT);
   G_1251GAT : And_gate port map( I1 => G_239GAT, I2 => G_477GAT, O => 
                           G_1251GAT_OUT);
   G_1248GAT : And_gate port map( I1 => G_239GAT, I2 => G_460GAT, O => 
                           G_1248GAT_OUT);
   G_1245GAT : And_gate port map( I1 => G_239GAT, I2 => G_443GAT, O => 
                           G_1245GAT_OUT);
   G_1242GAT : And_gate port map( I1 => G_239GAT, I2 => G_426GAT, O => 
                           G_1242GAT_OUT);
   G_1239GAT : And_gate port map( I1 => G_239GAT, I2 => G_409GAT, O => 
                           G_1239GAT_OUT);
   G_1236GAT : And_gate port map( I1 => G_239GAT, I2 => G_392GAT, O => 
                           G_1236GAT_OUT);
   G_1233GAT : And_gate port map( I1 => G_239GAT, I2 => G_375GAT, O => 
                           G_1233GAT_OUT);
   G_1230GAT : And_gate port map( I1 => G_239GAT, I2 => G_358GAT, O => 
                           G_1230GAT_OUT);
   G_1227GAT : And_gate port map( I1 => G_239GAT, I2 => G_341GAT, O => 
                           G_1227GAT_OUT);
   G_1224GAT : And_gate port map( I1 => G_239GAT, I2 => G_324GAT, O => 
                           G_1224GAT_OUT);
   G_1221GAT : And_gate port map( I1 => G_239GAT, I2 => G_307GAT, O => 
                           G_1221GAT_OUT);
   G_1218GAT : And_gate port map( I1 => G_239GAT, I2 => G_290GAT, O => 
                           G_1218GAT_OUT);
   G_1215GAT : And_gate port map( I1 => G_239GAT, I2 => G_273GAT, O => 
                           G_1215GAT_OUT);
   G_1212GAT : And_gate port map( I1 => G_222GAT, I2 => G_528GAT, O => 
                           G_1212GAT_OUT);
   G_1209GAT : And_gate port map( I1 => G_222GAT, I2 => G_511GAT, O => 
                           G_1209GAT_OUT);
   G_1206GAT : And_gate port map( I1 => G_222GAT, I2 => G_494GAT, O => 
                           G_1206GAT_OUT);
   G_1203GAT : And_gate port map( I1 => G_222GAT, I2 => G_477GAT, O => 
                           G_1203GAT_OUT);
   G_1200GAT : And_gate port map( I1 => G_222GAT, I2 => G_460GAT, O => 
                           G_1200GAT_OUT);
   G_1197GAT : And_gate port map( I1 => G_222GAT, I2 => G_443GAT, O => 
                           G_1197GAT_OUT);
   G_1194GAT : And_gate port map( I1 => G_222GAT, I2 => G_426GAT, O => 
                           G_1194GAT_OUT);
   G_1191GAT : And_gate port map( I1 => G_222GAT, I2 => G_409GAT, O => 
                           G_1191GAT_OUT);
   G_1188GAT : And_gate port map( I1 => G_222GAT, I2 => G_392GAT, O => 
                           G_1188GAT_OUT);
   G_1185GAT : And_gate port map( I1 => G_222GAT, I2 => G_375GAT, O => 
                           G_1185GAT_OUT);
   G_1182GAT : And_gate port map( I1 => G_222GAT, I2 => G_358GAT, O => 
                           G_1182GAT_OUT);
   G_1179GAT : And_gate port map( I1 => G_222GAT, I2 => G_341GAT, O => 
                           G_1179GAT_OUT);
   G_1176GAT : And_gate port map( I1 => G_222GAT, I2 => G_324GAT, O => 
                           G_1176GAT_OUT);
   G_1173GAT : And_gate port map( I1 => G_222GAT, I2 => G_307GAT, O => 
                           G_1173GAT_OUT);
   G_1170GAT : And_gate port map( I1 => G_222GAT, I2 => G_290GAT, O => 
                           G_1170GAT_OUT);
   G_1167GAT : And_gate port map( I1 => G_222GAT, I2 => G_273GAT, O => 
                           G_1167GAT_OUT);
   G_1164GAT : And_gate port map( I1 => G_205GAT, I2 => G_528GAT, O => 
                           G_1164GAT_OUT);
   G_1161GAT : And_gate port map( I1 => G_205GAT, I2 => G_511GAT, O => 
                           G_1161GAT_OUT);
   G_1158GAT : And_gate port map( I1 => G_205GAT, I2 => G_494GAT, O => 
                           G_1158GAT_OUT);
   G_1155GAT : And_gate port map( I1 => G_205GAT, I2 => G_477GAT, O => 
                           G_1155GAT_OUT);
   G_1152GAT : And_gate port map( I1 => G_205GAT, I2 => G_460GAT, O => 
                           G_1152GAT_OUT);
   G_1149GAT : And_gate port map( I1 => G_205GAT, I2 => G_443GAT, O => 
                           G_1149GAT_OUT);
   G_1146GAT : And_gate port map( I1 => G_205GAT, I2 => G_426GAT, O => 
                           G_1146GAT_OUT);
   G_1143GAT : And_gate port map( I1 => G_205GAT, I2 => G_409GAT, O => 
                           G_1143GAT_OUT);
   G_1140GAT : And_gate port map( I1 => G_205GAT, I2 => G_392GAT, O => 
                           G_1140GAT_OUT);
   G_1137GAT : And_gate port map( I1 => G_205GAT, I2 => G_375GAT, O => 
                           G_1137GAT_OUT);
   G_1134GAT : And_gate port map( I1 => G_205GAT, I2 => G_358GAT, O => 
                           G_1134GAT_OUT);
   G_1131GAT : And_gate port map( I1 => G_205GAT, I2 => G_341GAT, O => 
                           G_1131GAT_OUT);
   G_1128GAT : And_gate port map( I1 => G_205GAT, I2 => G_324GAT, O => 
                           G_1128GAT_OUT);
   G_1125GAT : And_gate port map( I1 => G_205GAT, I2 => G_307GAT, O => 
                           G_1125GAT_OUT);
   G_1122GAT : And_gate port map( I1 => G_205GAT, I2 => G_290GAT, O => 
                           G_1122GAT_OUT);
   G_1119GAT : And_gate port map( I1 => G_205GAT, I2 => G_273GAT, O => 
                           G_1119GAT_OUT);
   G_1116GAT : And_gate port map( I1 => G_188GAT, I2 => G_528GAT, O => 
                           G_1116GAT_OUT);
   G_1113GAT : And_gate port map( I1 => G_188GAT, I2 => G_511GAT, O => 
                           G_1113GAT_OUT);
   G_1110GAT : And_gate port map( I1 => G_188GAT, I2 => G_494GAT, O => 
                           G_1110GAT_OUT);
   G_1107GAT : And_gate port map( I1 => G_188GAT, I2 => G_477GAT, O => 
                           G_1107GAT_OUT);
   G_1104GAT : And_gate port map( I1 => G_188GAT, I2 => G_460GAT, O => 
                           G_1104GAT_OUT);
   G_1101GAT : And_gate port map( I1 => G_188GAT, I2 => G_443GAT, O => 
                           G_1101GAT_OUT);
   G_1098GAT : And_gate port map( I1 => G_188GAT, I2 => G_426GAT, O => 
                           G_1098GAT_OUT);
   G_1095GAT : And_gate port map( I1 => G_188GAT, I2 => G_409GAT, O => 
                           G_1095GAT_OUT);
   G_1092GAT : And_gate port map( I1 => G_188GAT, I2 => G_392GAT, O => 
                           G_1092GAT_OUT);
   G_1089GAT : And_gate port map( I1 => G_188GAT, I2 => G_375GAT, O => 
                           G_1089GAT_OUT);
   G_1086GAT : And_gate port map( I1 => G_188GAT, I2 => G_358GAT, O => 
                           G_1086GAT_OUT);
   G_1083GAT : And_gate port map( I1 => G_188GAT, I2 => G_341GAT, O => 
                           G_1083GAT_OUT);
   G_1080GAT : And_gate port map( I1 => G_188GAT, I2 => G_324GAT, O => 
                           G_1080GAT_OUT);
   G_1077GAT : And_gate port map( I1 => G_188GAT, I2 => G_307GAT, O => 
                           G_1077GAT_OUT);
   G_1074GAT : And_gate port map( I1 => G_188GAT, I2 => G_290GAT, O => 
                           G_1074GAT_OUT);
   G_1071GAT : And_gate port map( I1 => G_188GAT, I2 => G_273GAT, O => 
                           G_1071GAT_OUT);
   G_1068GAT : And_gate port map( I1 => G_171GAT, I2 => G_528GAT, O => 
                           G_1068GAT_OUT);
   G_1065GAT : And_gate port map( I1 => G_171GAT, I2 => G_511GAT, O => 
                           G_1065GAT_OUT);
   G_1062GAT : And_gate port map( I1 => G_171GAT, I2 => G_494GAT, O => 
                           G_1062GAT_OUT);
   G_1059GAT : And_gate port map( I1 => G_171GAT, I2 => G_477GAT, O => 
                           G_1059GAT_OUT);
   G_1056GAT : And_gate port map( I1 => G_171GAT, I2 => G_460GAT, O => 
                           G_1056GAT_OUT);
   G_1053GAT : And_gate port map( I1 => G_171GAT, I2 => G_443GAT, O => 
                           G_1053GAT_OUT);
   G_1050GAT : And_gate port map( I1 => G_171GAT, I2 => G_426GAT, O => 
                           G_1050GAT_OUT);
   G_1047GAT : And_gate port map( I1 => G_171GAT, I2 => G_409GAT, O => 
                           G_1047GAT_OUT);
   G_1044GAT : And_gate port map( I1 => G_171GAT, I2 => G_392GAT, O => 
                           G_1044GAT_OUT);
   G_1041GAT : And_gate port map( I1 => G_171GAT, I2 => G_375GAT, O => 
                           G_1041GAT_OUT);
   G_1038GAT : And_gate port map( I1 => G_171GAT, I2 => G_358GAT, O => 
                           G_1038GAT_OUT);
   G_1035GAT : And_gate port map( I1 => G_171GAT, I2 => G_341GAT, O => 
                           G_1035GAT_OUT);
   G_1032GAT : And_gate port map( I1 => G_171GAT, I2 => G_324GAT, O => 
                           G_1032GAT_OUT);
   G_1029GAT : And_gate port map( I1 => G_171GAT, I2 => G_307GAT, O => 
                           G_1029GAT_OUT);
   G_1026GAT : And_gate port map( I1 => G_171GAT, I2 => G_290GAT, O => 
                           G_1026GAT_OUT);
   G_1023GAT : And_gate port map( I1 => G_171GAT, I2 => G_273GAT, O => 
                           G_1023GAT_OUT);
   G_1020GAT : And_gate port map( I1 => G_154GAT, I2 => G_528GAT, O => 
                           G_1020GAT_OUT);
   G_1017GAT : And_gate port map( I1 => G_154GAT, I2 => G_511GAT, O => 
                           G_1017GAT_OUT);
   G_1014GAT : And_gate port map( I1 => G_154GAT, I2 => G_494GAT, O => 
                           G_1014GAT_OUT);
   G_1011GAT : And_gate port map( I1 => G_154GAT, I2 => G_477GAT, O => 
                           G_1011GAT_OUT);
   G_1008GAT : And_gate port map( I1 => G_154GAT, I2 => G_460GAT, O => 
                           G_1008GAT_OUT);
   G_1005GAT : And_gate port map( I1 => G_154GAT, I2 => G_443GAT, O => 
                           G_1005GAT_OUT);
   G_1002GAT : And_gate port map( I1 => G_154GAT, I2 => G_426GAT, O => 
                           G_1002GAT_OUT);
   G_999GAT : And_gate port map( I1 => G_154GAT, I2 => G_409GAT, O => 
                           G_999GAT_OUT);
   G_996GAT : And_gate port map( I1 => G_154GAT, I2 => G_392GAT, O => 
                           G_996GAT_OUT);
   G_993GAT : And_gate port map( I1 => G_154GAT, I2 => G_375GAT, O => 
                           G_993GAT_OUT);
   G_990GAT : And_gate port map( I1 => G_154GAT, I2 => G_358GAT, O => 
                           G_990GAT_OUT);
   G_987GAT : And_gate port map( I1 => G_154GAT, I2 => G_341GAT, O => 
                           G_987GAT_OUT);
   G_984GAT : And_gate port map( I1 => G_154GAT, I2 => G_324GAT, O => 
                           G_984GAT_OUT);
   G_981GAT : And_gate port map( I1 => G_154GAT, I2 => G_307GAT, O => 
                           G_981GAT_OUT);
   G_978GAT : And_gate port map( I1 => G_154GAT, I2 => G_290GAT, O => 
                           G_978GAT_OUT);
   G_975GAT : And_gate port map( I1 => G_154GAT, I2 => G_273GAT, O => 
                           G_975GAT_OUT);
   G_972GAT : And_gate port map( I1 => G_137GAT, I2 => G_528GAT, O => 
                           G_972GAT_OUT);
   G_969GAT : And_gate port map( I1 => G_137GAT, I2 => G_511GAT, O => 
                           G_969GAT_OUT);
   G_966GAT : And_gate port map( I1 => G_137GAT, I2 => G_494GAT, O => 
                           G_966GAT_OUT);
   G_963GAT : And_gate port map( I1 => G_137GAT, I2 => G_477GAT, O => 
                           G_963GAT_OUT);
   G_960GAT : And_gate port map( I1 => G_137GAT, I2 => G_460GAT, O => 
                           G_960GAT_OUT);
   G_957GAT : And_gate port map( I1 => G_137GAT, I2 => G_443GAT, O => 
                           G_957GAT_OUT);
   G_954GAT : And_gate port map( I1 => G_137GAT, I2 => G_426GAT, O => 
                           G_954GAT_OUT);
   G_951GAT : And_gate port map( I1 => G_137GAT, I2 => G_409GAT, O => 
                           G_951GAT_OUT);
   G_948GAT : And_gate port map( I1 => G_137GAT, I2 => G_392GAT, O => 
                           G_948GAT_OUT);
   G_945GAT : And_gate port map( I1 => G_137GAT, I2 => G_375GAT, O => 
                           G_945GAT_OUT);
   G_942GAT : And_gate port map( I1 => G_137GAT, I2 => G_358GAT, O => 
                           G_942GAT_OUT);
   G_939GAT : And_gate port map( I1 => G_137GAT, I2 => G_341GAT, O => 
                           G_939GAT_OUT);
   G_936GAT : And_gate port map( I1 => G_137GAT, I2 => G_324GAT, O => 
                           G_936GAT_OUT);
   G_933GAT : And_gate port map( I1 => G_137GAT, I2 => G_307GAT, O => 
                           G_933GAT_OUT);
   G_930GAT : And_gate port map( I1 => G_137GAT, I2 => G_290GAT, O => 
                           G_930GAT_OUT);
   G_927GAT : And_gate port map( I1 => G_137GAT, I2 => G_273GAT, O => 
                           G_927GAT_OUT);
   G_924GAT : And_gate port map( I1 => G_120GAT, I2 => G_528GAT, O => 
                           G_924GAT_OUT);
   G_921GAT : And_gate port map( I1 => G_120GAT, I2 => G_511GAT, O => 
                           G_921GAT_OUT);
   G_918GAT : And_gate port map( I1 => G_120GAT, I2 => G_494GAT, O => 
                           G_918GAT_OUT);
   G_915GAT : And_gate port map( I1 => G_120GAT, I2 => G_477GAT, O => 
                           G_915GAT_OUT);
   G_912GAT : And_gate port map( I1 => G_120GAT, I2 => G_460GAT, O => 
                           G_912GAT_OUT);
   G_909GAT : And_gate port map( I1 => G_120GAT, I2 => G_443GAT, O => 
                           G_909GAT_OUT);
   G_906GAT : And_gate port map( I1 => G_120GAT, I2 => G_426GAT, O => 
                           G_906GAT_OUT);
   G_903GAT : And_gate port map( I1 => G_120GAT, I2 => G_409GAT, O => 
                           G_903GAT_OUT);
   G_900GAT : And_gate port map( I1 => G_120GAT, I2 => G_392GAT, O => 
                           G_900GAT_OUT);
   G_897GAT : And_gate port map( I1 => G_120GAT, I2 => G_375GAT, O => 
                           G_897GAT_OUT);
   G_894GAT : And_gate port map( I1 => G_120GAT, I2 => G_358GAT, O => 
                           G_894GAT_OUT);
   G_891GAT : And_gate port map( I1 => G_120GAT, I2 => G_341GAT, O => 
                           G_891GAT_OUT);
   G_888GAT : And_gate port map( I1 => G_120GAT, I2 => G_324GAT, O => 
                           G_888GAT_OUT);
   G_885GAT : And_gate port map( I1 => G_120GAT, I2 => G_307GAT, O => 
                           G_885GAT_OUT);
   G_882GAT : And_gate port map( I1 => G_120GAT, I2 => G_290GAT, O => 
                           G_882GAT_OUT);
   G_879GAT : And_gate port map( I1 => G_120GAT, I2 => G_273GAT, O => 
                           G_879GAT_OUT);
   G_876GAT : And_gate port map( I1 => G_103GAT, I2 => G_528GAT, O => 
                           G_876GAT_OUT);
   G_873GAT : And_gate port map( I1 => G_103GAT, I2 => G_511GAT, O => 
                           G_873GAT_OUT);
   G_870GAT : And_gate port map( I1 => G_103GAT, I2 => G_494GAT, O => 
                           G_870GAT_OUT);
   G_867GAT : And_gate port map( I1 => G_103GAT, I2 => G_477GAT, O => 
                           G_867GAT_OUT);
   G_864GAT : And_gate port map( I1 => G_103GAT, I2 => G_460GAT, O => 
                           G_864GAT_OUT);
   G_861GAT : And_gate port map( I1 => G_103GAT, I2 => G_443GAT, O => 
                           G_861GAT_OUT);
   G_858GAT : And_gate port map( I1 => G_103GAT, I2 => G_426GAT, O => 
                           G_858GAT_OUT);
   G_855GAT : And_gate port map( I1 => G_103GAT, I2 => G_409GAT, O => 
                           G_855GAT_OUT);
   G_852GAT : And_gate port map( I1 => G_103GAT, I2 => G_392GAT, O => 
                           G_852GAT_OUT);
   G_849GAT : And_gate port map( I1 => G_103GAT, I2 => G_375GAT, O => 
                           G_849GAT_OUT);
   G_846GAT : And_gate port map( I1 => G_103GAT, I2 => G_358GAT, O => 
                           G_846GAT_OUT);
   G_843GAT : And_gate port map( I1 => G_103GAT, I2 => G_341GAT, O => 
                           G_843GAT_OUT);
   G_840GAT : And_gate port map( I1 => G_103GAT, I2 => G_324GAT, O => 
                           G_840GAT_OUT);
   G_837GAT : And_gate port map( I1 => G_103GAT, I2 => G_307GAT, O => 
                           G_837GAT_OUT);
   G_834GAT : And_gate port map( I1 => G_103GAT, I2 => G_290GAT, O => 
                           G_834GAT_OUT);
   G_831GAT : And_gate port map( I1 => G_103GAT, I2 => G_273GAT, O => 
                           G_831GAT_OUT);
   G_828GAT : And_gate port map( I1 => G_86GAT, I2 => G_528GAT, O => 
                           G_828GAT_OUT);
   G_825GAT : And_gate port map( I1 => G_86GAT, I2 => G_511GAT, O => 
                           G_825GAT_OUT);
   G_822GAT : And_gate port map( I1 => G_86GAT, I2 => G_494GAT, O => 
                           G_822GAT_OUT);
   G_819GAT : And_gate port map( I1 => G_86GAT, I2 => G_477GAT, O => 
                           G_819GAT_OUT);
   G_816GAT : And_gate port map( I1 => G_86GAT, I2 => G_460GAT, O => 
                           G_816GAT_OUT);
   G_813GAT : And_gate port map( I1 => G_86GAT, I2 => G_443GAT, O => 
                           G_813GAT_OUT);
   G_810GAT : And_gate port map( I1 => G_86GAT, I2 => G_426GAT, O => 
                           G_810GAT_OUT);
   G_807GAT : And_gate port map( I1 => G_86GAT, I2 => G_409GAT, O => 
                           G_807GAT_OUT);
   G_804GAT : And_gate port map( I1 => G_86GAT, I2 => G_392GAT, O => 
                           G_804GAT_OUT);
   G_801GAT : And_gate port map( I1 => G_86GAT, I2 => G_375GAT, O => 
                           G_801GAT_OUT);
   G_798GAT : And_gate port map( I1 => G_86GAT, I2 => G_358GAT, O => 
                           G_798GAT_OUT);
   G_795GAT : And_gate port map( I1 => G_86GAT, I2 => G_341GAT, O => 
                           G_795GAT_OUT);
   G_792GAT : And_gate port map( I1 => G_86GAT, I2 => G_324GAT, O => 
                           G_792GAT_OUT);
   G_789GAT : And_gate port map( I1 => G_86GAT, I2 => G_307GAT, O => 
                           G_789GAT_OUT);
   G_786GAT : And_gate port map( I1 => G_86GAT, I2 => G_290GAT, O => 
                           G_786GAT_OUT);
   G_783GAT : And_gate port map( I1 => G_86GAT, I2 => G_273GAT, O => 
                           G_783GAT_OUT);
   G_780GAT : And_gate port map( I1 => G_69GAT, I2 => G_528GAT, O => 
                           G_780GAT_OUT);
   G_777GAT : And_gate port map( I1 => G_69GAT, I2 => G_511GAT, O => 
                           G_777GAT_OUT);
   G_774GAT : And_gate port map( I1 => G_69GAT, I2 => G_494GAT, O => 
                           G_774GAT_OUT);
   G_771GAT : And_gate port map( I1 => G_69GAT, I2 => G_477GAT, O => 
                           G_771GAT_OUT);
   G_768GAT : And_gate port map( I1 => G_69GAT, I2 => G_460GAT, O => 
                           G_768GAT_OUT);
   G_765GAT : And_gate port map( I1 => G_69GAT, I2 => G_443GAT, O => 
                           G_765GAT_OUT);
   G_762GAT : And_gate port map( I1 => G_69GAT, I2 => G_426GAT, O => 
                           G_762GAT_OUT);
   G_759GAT : And_gate port map( I1 => G_69GAT, I2 => G_409GAT, O => 
                           G_759GAT_OUT);
   G_756GAT : And_gate port map( I1 => G_69GAT, I2 => G_392GAT, O => 
                           G_756GAT_OUT);
   G_753GAT : And_gate port map( I1 => G_69GAT, I2 => G_375GAT, O => 
                           G_753GAT_OUT);
   G_750GAT : And_gate port map( I1 => G_69GAT, I2 => G_358GAT, O => 
                           G_750GAT_OUT);
   G_747GAT : And_gate port map( I1 => G_69GAT, I2 => G_341GAT, O => 
                           G_747GAT_OUT);
   G_744GAT : And_gate port map( I1 => G_69GAT, I2 => G_324GAT, O => 
                           G_744GAT_OUT);
   G_741GAT : And_gate port map( I1 => G_69GAT, I2 => G_307GAT, O => 
                           G_741GAT_OUT);
   G_738GAT : And_gate port map( I1 => G_69GAT, I2 => G_290GAT, O => 
                           G_738GAT_OUT);
   G_735GAT : And_gate port map( I1 => G_69GAT, I2 => G_273GAT, O => 
                           G_735GAT_OUT);
   G_732GAT : And_gate port map( I1 => G_52GAT, I2 => G_528GAT, O => 
                           G_732GAT_OUT);
   G_729GAT : And_gate port map( I1 => G_52GAT, I2 => G_511GAT, O => 
                           G_729GAT_OUT);
   G_726GAT : And_gate port map( I1 => G_52GAT, I2 => G_494GAT, O => 
                           G_726GAT_OUT);
   G_723GAT : And_gate port map( I1 => G_52GAT, I2 => G_477GAT, O => 
                           G_723GAT_OUT);
   G_720GAT : And_gate port map( I1 => G_52GAT, I2 => G_460GAT, O => 
                           G_720GAT_OUT);
   G_717GAT : And_gate port map( I1 => G_52GAT, I2 => G_443GAT, O => 
                           G_717GAT_OUT);
   G_714GAT : And_gate port map( I1 => G_52GAT, I2 => G_426GAT, O => 
                           G_714GAT_OUT);
   G_711GAT : And_gate port map( I1 => G_52GAT, I2 => G_409GAT, O => 
                           G_711GAT_OUT);
   G_708GAT : And_gate port map( I1 => G_52GAT, I2 => G_392GAT, O => 
                           G_708GAT_OUT);
   G_705GAT : And_gate port map( I1 => G_52GAT, I2 => G_375GAT, O => 
                           G_705GAT_OUT);
   G_702GAT : And_gate port map( I1 => G_52GAT, I2 => G_358GAT, O => 
                           G_702GAT_OUT);
   G_699GAT : And_gate port map( I1 => G_52GAT, I2 => G_341GAT, O => 
                           G_699GAT_OUT);
   G_696GAT : And_gate port map( I1 => G_52GAT, I2 => G_324GAT, O => 
                           G_696GAT_OUT);
   G_693GAT : And_gate port map( I1 => G_52GAT, I2 => G_307GAT, O => 
                           G_693GAT_OUT);
   G_690GAT : And_gate port map( I1 => G_52GAT, I2 => G_290GAT, O => 
                           G_690GAT_OUT);
   G_687GAT : And_gate port map( I1 => G_52GAT, I2 => G_273GAT, O => 
                           G_687GAT_OUT);
   G_684GAT : And_gate port map( I1 => G_35GAT, I2 => G_528GAT, O => 
                           G_684GAT_OUT);
   G_681GAT : And_gate port map( I1 => G_35GAT, I2 => G_511GAT, O => 
                           G_681GAT_OUT);
   G_678GAT : And_gate port map( I1 => G_35GAT, I2 => G_494GAT, O => 
                           G_678GAT_OUT);
   G_675GAT : And_gate port map( I1 => G_35GAT, I2 => G_477GAT, O => 
                           G_675GAT_OUT);
   G_672GAT : And_gate port map( I1 => G_35GAT, I2 => G_460GAT, O => 
                           G_672GAT_OUT);
   G_669GAT : And_gate port map( I1 => G_35GAT, I2 => G_443GAT, O => 
                           G_669GAT_OUT);
   G_666GAT : And_gate port map( I1 => G_35GAT, I2 => G_426GAT, O => 
                           G_666GAT_OUT);
   G_663GAT : And_gate port map( I1 => G_35GAT, I2 => G_409GAT, O => 
                           G_663GAT_OUT);
   G_660GAT : And_gate port map( I1 => G_35GAT, I2 => G_392GAT, O => 
                           G_660GAT_OUT);
   G_657GAT : And_gate port map( I1 => G_35GAT, I2 => G_375GAT, O => 
                           G_657GAT_OUT);
   G_654GAT : And_gate port map( I1 => G_35GAT, I2 => G_358GAT, O => 
                           G_654GAT_OUT);
   G_651GAT : And_gate port map( I1 => G_35GAT, I2 => G_341GAT, O => 
                           G_651GAT_OUT);
   G_648GAT : And_gate port map( I1 => G_35GAT, I2 => G_324GAT, O => 
                           G_648GAT_OUT);
   G_645GAT : And_gate port map( I1 => G_35GAT, I2 => G_307GAT, O => 
                           G_645GAT_OUT);
   G_642GAT : And_gate port map( I1 => G_35GAT, I2 => G_290GAT, O => 
                           G_642GAT_OUT);
   G_639GAT : And_gate port map( I1 => G_35GAT, I2 => G_273GAT, O => 
                           G_639GAT_OUT);
   G_636GAT : And_gate port map( I1 => G_18GAT, I2 => G_528GAT, O => 
                           G_636GAT_OUT);
   G_633GAT : And_gate port map( I1 => G_18GAT, I2 => G_511GAT, O => 
                           G_633GAT_OUT);
   G_630GAT : And_gate port map( I1 => G_18GAT, I2 => G_494GAT, O => 
                           G_630GAT_OUT);
   G_627GAT : And_gate port map( I1 => G_18GAT, I2 => G_477GAT, O => 
                           G_627GAT_OUT);
   G_624GAT : And_gate port map( I1 => G_18GAT, I2 => G_460GAT, O => 
                           G_624GAT_OUT);
   G_621GAT : And_gate port map( I1 => G_18GAT, I2 => G_443GAT, O => 
                           G_621GAT_OUT);
   G_618GAT : And_gate port map( I1 => G_18GAT, I2 => G_426GAT, O => 
                           G_618GAT_OUT);
   G_615GAT : And_gate port map( I1 => G_18GAT, I2 => G_409GAT, O => 
                           G_615GAT_OUT);
   G_612GAT : And_gate port map( I1 => G_18GAT, I2 => G_392GAT, O => 
                           G_612GAT_OUT);
   G_609GAT : And_gate port map( I1 => G_18GAT, I2 => G_375GAT, O => 
                           G_609GAT_OUT);
   G_606GAT : And_gate port map( I1 => G_18GAT, I2 => G_358GAT, O => 
                           G_606GAT_OUT);
   G_603GAT : And_gate port map( I1 => G_18GAT, I2 => G_341GAT, O => 
                           G_603GAT_OUT);
   G_600GAT : And_gate port map( I1 => G_18GAT, I2 => G_324GAT, O => 
                           G_600GAT_OUT);
   G_597GAT : And_gate port map( I1 => G_18GAT, I2 => G_307GAT, O => 
                           G_597GAT_OUT);
   G_594GAT : And_gate port map( I1 => G_18GAT, I2 => G_290GAT, O => 
                           G_594GAT_OUT);
   G_591GAT : And_gate port map( I1 => G_18GAT, I2 => G_273GAT, O => 
                           G_591GAT_OUT);
   G_588GAT : And_gate port map( I1 => G_1GAT, I2 => G_528GAT, O => 
                           G_588GAT_OUT);
   G_585GAT : And_gate port map( I1 => G_1GAT, I2 => G_511GAT, O => 
                           G_585GAT_OUT);
   G_582GAT : And_gate port map( I1 => G_1GAT, I2 => G_494GAT, O => 
                           G_582GAT_OUT);
   G_579GAT : And_gate port map( I1 => G_1GAT, I2 => G_477GAT, O => 
                           G_579GAT_OUT);
   G_576GAT : And_gate port map( I1 => G_1GAT, I2 => G_460GAT, O => 
                           G_576GAT_OUT);
   G_573GAT : And_gate port map( I1 => G_1GAT, I2 => G_443GAT, O => 
                           G_573GAT_OUT);
   G_570GAT : And_gate port map( I1 => G_1GAT, I2 => G_426GAT, O => 
                           G_570GAT_OUT);
   G_567GAT : And_gate port map( I1 => G_1GAT, I2 => G_409GAT, O => 
                           G_567GAT_OUT);
   G_564GAT : And_gate port map( I1 => G_1GAT, I2 => G_392GAT, O => 
                           G_564GAT_OUT);
   G_561GAT : And_gate port map( I1 => G_1GAT, I2 => G_375GAT, O => 
                           G_561GAT_OUT);
   G_558GAT : And_gate port map( I1 => G_1GAT, I2 => G_358GAT, O => 
                           G_558GAT_OUT);
   G_555GAT : And_gate port map( I1 => G_1GAT, I2 => G_341GAT, O => 
                           G_555GAT_OUT);
   G_552GAT : And_gate port map( I1 => G_1GAT, I2 => G_324GAT, O => 
                           G_552GAT_OUT);
   G_549GAT : And_gate port map( I1 => G_1GAT, I2 => G_307GAT, O => 
                           G_549GAT_OUT);
   G_546GAT : And_gate port map( I1 => G_1GAT, I2 => G_290GAT, O => 
                           G_546GAT_OUT);
   G_545GAT : And_gate port map( I1 => G_1GAT, I2 => G_273GAT, O => G_545GAT_PO
                           );
   G_1581GAT : Nor_gate port map( I1 => G_1506GAT_OUT, I2 => G_1507GAT_OUT, O 
                           => G_1581GAT_PO);
   G_1901GAT : Nor_gate port map( I1 => G_1824GAT_OUT, I2 => G_1825GAT_OUT, O 
                           => G_1901GAT_PO);
   G_2223GAT : Nor_gate port map( I1 => G_2149GAT_OUT, I2 => G_2150GAT_OUT, O 
                           => G_2223GAT_PO);
   G_2548GAT : Nor_gate port map( I1 => G_2476GAT_OUT, I2 => G_2477GAT_OUT, O 
                           => G_2548GAT_PO);
   G_2877GAT : Nor_gate port map( I1 => G_2806GAT_OUT, I2 => G_2807GAT_OUT, O 
                           => G_2877GAT_PO);
   G_3211GAT : Nor_gate port map( I1 => G_3140GAT_OUT, I2 => G_3141GAT_OUT, O 
                           => G_3211GAT_PO);
   G_3552GAT : Nor_gate port map( I1 => G_3479GAT_OUT, I2 => G_3480GAT_OUT, O 
                           => G_3552GAT_PO);
   G_3895GAT : Nor_gate port map( I1 => G_3825GAT_OUT, I2 => G_3826GAT_OUT, O 
                           => G_3895GAT_PO);
   G_4241GAT : Nor_gate port map( I1 => G_4173GAT_OUT, I2 => G_4174GAT_OUT, O 
                           => G_4241GAT_PO);
   G_4591GAT : Nor_gate port map( I1 => G_4524GAT_OUT, I2 => G_4525GAT_OUT, O 
                           => G_4591GAT_PO);
   G_4946GAT : Nor_gate port map( I1 => G_4879GAT_OUT, I2 => G_4880GAT_OUT, O 
                           => G_4946GAT_PO);
   G_5308GAT : Nor_gate port map( I1 => G_5239GAT_OUT, I2 => G_5240GAT_OUT, O 
                           => G_5308GAT_PO);
   G_5672GAT : Nor_gate port map( I1 => G_5606GAT_OUT, I2 => G_5607GAT_OUT, O 
                           => G_5672GAT_PO);
   G_5971GAT : Nor_gate port map( I1 => G_5928GAT_OUT, I2 => G_5929GAT_OUT, O 
                           => G_5971GAT_PO);
   G_6123GAT : Nor_gate port map( I1 => G_6106GAT_OUT, I2 => G_6107GAT_OUT, O 
                           => G_6123GAT_PO);
   G_6150GAT : Nor_gate port map( I1 => G_6145GAT_OUT, I2 => G_6146GAT_OUT, O 
                           => G_6150GAT_PO);
   G_6160GAT : Nor_gate port map( I1 => G_6155GAT_OUT, I2 => G_6156GAT_OUT, O 
                           => G_6160GAT_PO);
   G_6170GAT : Nor_gate port map( I1 => G_6165GAT_OUT, I2 => G_6166GAT_OUT, O 
                           => G_6170GAT_PO);
   G_6180GAT : Nor_gate port map( I1 => G_6175GAT_OUT, I2 => G_6176GAT_OUT, O 
                           => G_6180GAT_PO);
   G_6190GAT : Nor_gate port map( I1 => G_6185GAT_OUT, I2 => G_6186GAT_OUT, O 
                           => G_6190GAT_PO);
   G_6200GAT : Nor_gate port map( I1 => G_6195GAT_OUT, I2 => G_6196GAT_OUT, O 
                           => G_6200GAT_PO);
   G_6210GAT : Nor_gate port map( I1 => G_6205GAT_OUT, I2 => G_6206GAT_OUT, O 
                           => G_6210GAT_PO);
   G_6220GAT : Nor_gate port map( I1 => G_6215GAT_OUT, I2 => G_6216GAT_OUT, O 
                           => G_6220GAT_PO);
   G_6230GAT : Nor_gate port map( I1 => G_6225GAT_OUT, I2 => G_6226GAT_OUT, O 
                           => G_6230GAT_PO);
   G_6240GAT : Nor_gate port map( I1 => G_6235GAT_OUT, I2 => G_6236GAT_OUT, O 
                           => G_6240GAT_PO);
   G_6250GAT : Nor_gate port map( I1 => G_6245GAT_OUT, I2 => G_6246GAT_OUT, O 
                           => G_6250GAT_PO);
   G_6260GAT : Nor_gate port map( I1 => G_6255GAT_OUT, I2 => G_6256GAT_OUT, O 
                           => G_6260GAT_PO);
   G_6270GAT : Nor_gate port map( I1 => G_6265GAT_OUT, I2 => G_6266GAT_OUT, O 
                           => G_6270GAT_PO);
   G_6280GAT : Nor_gate port map( I1 => G_6275GAT_OUT, I2 => G_6276GAT_OUT, O 
                           => G_6280GAT_PO);
   G_6287GAT : Nor_gate port map( I1 => G_5602GAT_OUT, I2 => G_6281GAT_OUT, O 
                           => G_6287GAT_PO);
   G_6288GAT : Nor_gate port map( I1 => G_6285GAT_OUT, I2 => G_6286GAT_OUT, O 
                           => G_6288GAT_PO);

end SYN_USE_DEFA_ARCH_NAME;
